`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module rvdm( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [1:0]  io_dmi_req_bits_op, // @[:@6.4]
  input  [6:0]  io_dmi_req_bits_addr, // @[:@6.4]
  input  [31:0] io_dmi_req_bits_data, // @[:@6.4]
  input         io_dmi_req_valid, // @[:@6.4]
  output        io_dmi_req_ready, // @[:@6.4]
  output [1:0]  io_dmi_resp_bits_resp, // @[:@6.4]
  output [31:0] io_dmi_resp_bits_data, // @[:@6.4]
  output        io_dmi_resp_valid, // @[:@6.4]
  output [4:0]  io_ddpath_addr, // @[:@6.4]
  output [31:0] io_ddpath_wdata, // @[:@6.4]
  output        io_ddpath_valid, // @[:@6.4]
  input  [31:0] io_ddpath_rdata, // @[:@6.4]
  output [31:0] io_ddmem_req_addr, // @[:@6.4]
  output [31:0] io_ddmem_req_data, // @[:@6.4]
  output        io_ddmem_req_mfunc, // @[:@6.4]
  output        io_ddmem_req_valid, // @[:@6.4]
  input         io_ddmem_req_ready, // @[:@6.4]
  input  [31:0] io_ddmem_resp_data, // @[:@6.4]
  input         io_ddmem_resp_valid, // @[:@6.4]
  output        io_rstcore // @[:@6.4]
);
  reg [31:0] reg_dmstatus; // @[rvdm.scala 219:27:@32.4]
  reg [31:0] _RAND_0;
  reg [31:0] reg_dmcontrol; // @[rvdm.scala 220:28:@33.4]
  reg [31:0] _RAND_1;
  reg [31:0] reg_sbcs; // @[rvdm.scala 221:23:@34.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_abstractcs; // @[rvdm.scala 222:29:@35.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_command; // @[rvdm.scala 223:26:@36.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_progbuf_0; // @[rvdm.scala 224:26:@37.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_data_0; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_data_1; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_7;
  reg [31:0] reg_data_2; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_8;
  reg [31:0] reg_data_3; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_9;
  reg [31:0] reg_data_4; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_10;
  reg [31:0] reg_data_5; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_11;
  reg [31:0] reg_data_6; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_12;
  reg [31:0] reg_data_7; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_13;
  reg [31:0] reg_data_8; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_14;
  reg [31:0] reg_data_9; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_15;
  reg [31:0] reg_data_10; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_16;
  reg [31:0] reg_data_11; // @[rvdm.scala 225:23:@38.4]
  reg [31:0] _RAND_17;
  reg [31:0] reg_sbaddress_0; // @[rvdm.scala 227:28:@39.4]
  reg [31:0] _RAND_18;
  reg [31:0] reg_sbaddress_1; // @[rvdm.scala 227:28:@39.4]
  reg [31:0] _RAND_19;
  reg [31:0] reg_sbaddress_2; // @[rvdm.scala 227:28:@39.4]
  reg [31:0] _RAND_20;
  reg [31:0] reg_sbdata_0; // @[rvdm.scala 228:25:@40.4]
  reg [31:0] _RAND_21;
  reg  reg_regrw; // @[rvdm.scala 230:24:@41.4]
  reg [31:0] _RAND_22;
  reg  reg_mrdata_requested; // @[rvdm.scala 233:35:@42.4]
  reg [31:0] _RAND_23;
  reg  reg_delay_mrwdata_valid; // @[rvdm.scala 234:38:@43.4]
  reg [31:0] _RAND_24;
  reg  reg_ddmem_req_valid; // @[rvdm.scala 236:34:@44.4]
  reg [31:0] _RAND_25;
  reg  reg_rstcore; // @[rvdm.scala 238:26:@45.4]
  reg [31:0] _RAND_26;
  wire  _T_132; // @[rvdm.scala 278:74:@51.4]
  wire  _T_144; // @[rvdm.scala 278:74:@57.4]
  wire  _T_146; // @[rvdm.scala 278:74:@58.4]
  wire  _T_154; // @[rvdm.scala 278:74:@62.4]
  wire  _T_156; // @[rvdm.scala 278:74:@63.4]
  wire  _T_158; // @[rvdm.scala 278:74:@64.4]
  wire  _T_160; // @[rvdm.scala 278:74:@65.4]
  wire  _T_162; // @[rvdm.scala 278:74:@66.4]
  wire  _T_164; // @[rvdm.scala 278:74:@67.4]
  wire  _T_166; // @[rvdm.scala 278:74:@68.4]
  wire  _T_168; // @[rvdm.scala 278:74:@69.4]
  wire  _T_170; // @[rvdm.scala 278:74:@70.4]
  wire  _T_172; // @[rvdm.scala 278:74:@71.4]
  wire  _T_174; // @[rvdm.scala 278:74:@72.4]
  wire  _T_176; // @[rvdm.scala 278:74:@73.4]
  wire  _T_178; // @[rvdm.scala 278:74:@74.4]
  wire  _T_212; // @[rvdm.scala 278:74:@91.4]
  wire  _T_214; // @[rvdm.scala 278:74:@92.4]
  wire  _T_216; // @[rvdm.scala 278:74:@93.4]
  wire  _T_218; // @[rvdm.scala 278:74:@94.4]
  wire [29:0] _T_277; // @[:@100.4]
  wire [3:0] _T_278; // @[rvdm.scala 290:42:@102.4]
  wire  dmstatus_devtreevalid; // @[rvdm.scala 290:42:@104.4]
  wire  dmstatus_rsrvd4; // @[rvdm.scala 290:42:@106.4]
  wire  dmstatus_authbusy; // @[rvdm.scala 290:42:@108.4]
  wire  _T_282; // @[rvdm.scala 290:42:@110.4]
  wire  dmstatus_anyhalted; // @[rvdm.scala 290:42:@112.4]
  wire  dmstatus_anyrunning; // @[rvdm.scala 290:42:@116.4]
  wire  dmstatus_anyunavail; // @[rvdm.scala 290:42:@120.4]
  wire  dmstatus_allunavail; // @[rvdm.scala 290:42:@122.4]
  wire  dmstatus_anynonexistent; // @[rvdm.scala 290:42:@124.4]
  wire  dmstatus_allnonexistent; // @[rvdm.scala 290:42:@126.4]
  wire  dmstatus_allresumeack; // @[rvdm.scala 290:42:@128.4]
  wire  dmstatus_anyhavereset; // @[rvdm.scala 290:42:@130.4]
  wire  dmstatus_allhavereset; // @[rvdm.scala 290:42:@132.4]
  wire  dmstatus_rsrvd3; // @[rvdm.scala 290:42:@134.4]
  wire  dmstatus_impebreak; // @[rvdm.scala 290:42:@136.4]
  wire  dmstatus_rsrvd2; // @[rvdm.scala 290:42:@138.4]
  wire [2:0] dmstatus_dmerr; // @[rvdm.scala 290:42:@140.4]
  wire [4:0] dmstatus_rsrvd1; // @[rvdm.scala 290:42:@142.4]
  wire  _T_305; // @[rvdm.scala 292:44:@169.4]
  wire  _T_306; // @[rvdm.scala 292:44:@171.4]
  wire [13:0] dmcontrol_rsrvd2; // @[rvdm.scala 292:44:@173.4]
  wire [9:0] dmcontrol_hartsel; // @[rvdm.scala 292:44:@175.4]
  wire  dmcontrol_hasel; // @[rvdm.scala 292:44:@177.4]
  wire  dmcontrol_rsrvd1; // @[rvdm.scala 292:44:@179.4]
  wire  dmcontrol_ackharvereset; // @[rvdm.scala 292:44:@181.4]
  wire  _T_312; // @[rvdm.scala 292:44:@183.4]
  wire  _T_313; // @[rvdm.scala 292:44:@185.4]
  wire  _T_314; // @[rvdm.scala 292:44:@187.4]
  wire  sbcs_sbaccess8; // @[rvdm.scala 294:34:@203.4]
  wire  sbcs_sbaccess16; // @[rvdm.scala 294:34:@205.4]
  wire  _T_323; // @[rvdm.scala 294:34:@207.4]
  wire  sbcs_sbaccess64; // @[rvdm.scala 294:34:@209.4]
  wire  sbcs_sbaccess128; // @[rvdm.scala 294:34:@211.4]
  wire [6:0] _T_326; // @[rvdm.scala 294:34:@213.4]
  wire [2:0] _T_327; // @[rvdm.scala 294:34:@215.4]
  wire  _T_328; // @[rvdm.scala 294:34:@217.4]
  wire  _T_329; // @[rvdm.scala 294:34:@219.4]
  wire [2:0] _T_330; // @[rvdm.scala 294:34:@221.4]
  wire  _T_331; // @[rvdm.scala 294:34:@223.4]
  wire [10:0] sbcs_rsrvd1; // @[rvdm.scala 294:34:@225.4]
  wire [4:0] _T_339; // @[rvdm.scala 296:46:@243.4]
  wire [2:0] abstractcs_rsrvd4; // @[rvdm.scala 296:46:@245.4]
  wire [2:0] _T_341; // @[rvdm.scala 296:46:@247.4]
  wire  abstractcs_rsrvd3; // @[rvdm.scala 296:46:@249.4]
  wire  abstractcs_busy; // @[rvdm.scala 296:46:@251.4]
  wire [10:0] abstractcs_rsrvd2; // @[rvdm.scala 296:46:@253.4]
  wire [4:0] _T_345; // @[rvdm.scala 296:46:@255.4]
  wire [2:0] abstractcs_rsrvd1; // @[rvdm.scala 296:46:@257.4]
  wire [15:0] _T_353; // @[rvdm.scala 298:40:@271.4]
  wire  _T_354; // @[rvdm.scala 298:40:@273.4]
  wire  _T_355; // @[rvdm.scala 298:40:@275.4]
  wire  _T_356; // @[rvdm.scala 298:40:@277.4]
  wire  command_rsrvd2; // @[rvdm.scala 298:40:@279.4]
  wire [2:0] command_size; // @[rvdm.scala 298:40:@281.4]
  wire  command_rsrvd1; // @[rvdm.scala 298:40:@283.4]
  wire [7:0] command_cmdtype; // @[rvdm.scala 298:40:@285.4]
  wire [3:0] dmstatus_version; // @[rvdm.scala 498:26:@735.4]
  wire [4:0] _T_361; // @[rvdm.scala 302:30:@297.4]
  wire  dmstatus_authenticated; // @[rvdm.scala 498:26:@735.4]
  wire [1:0] _T_362; // @[rvdm.scala 302:30:@298.4]
  wire [2:0] _T_363; // @[rvdm.scala 302:30:@299.4]
  wire [7:0] _T_364; // @[rvdm.scala 302:30:@300.4]
  wire  _T_384; // @[rvdm.scala 306:29:@321.4]
  wire  _T_461; // @[rvdm.scala 342:59:@441.8]
  wire  _GEN_22; // @[rvdm.scala 341:42:@419.6]
  wire  dmcontrol_haltreq; // @[rvdm.scala 306:50:@322.4]
  wire [1:0] _T_365; // @[rvdm.scala 302:30:@301.4]
  wire  _T_460; // @[rvdm.scala 342:59:@439.8]
  wire  _GEN_23; // @[rvdm.scala 341:42:@419.6]
  wire  dmcontrol_resumereq; // @[rvdm.scala 306:50:@322.4]
  wire [1:0] _T_366; // @[rvdm.scala 302:30:@302.4]
  wire [2:0] _T_367; // @[rvdm.scala 302:30:@303.4]
  wire [4:0] _T_368; // @[rvdm.scala 302:30:@304.4]
  wire [12:0] _T_369; // @[rvdm.scala 302:30:@305.4]
  wire [1:0] _T_370; // @[rvdm.scala 302:30:@306.4]
  wire [1:0] _T_371; // @[rvdm.scala 302:30:@307.4]
  wire [2:0] _T_372; // @[rvdm.scala 302:30:@308.4]
  wire [4:0] _T_373; // @[rvdm.scala 302:30:@309.4]
  wire [1:0] _T_374; // @[rvdm.scala 302:30:@310.4]
  wire [2:0] _T_375; // @[rvdm.scala 302:30:@311.4]
  wire [7:0] _T_376; // @[rvdm.scala 302:30:@312.4]
  wire [8:0] _T_377; // @[rvdm.scala 302:30:@313.4]
  wire [11:0] _T_378; // @[rvdm.scala 302:30:@314.4]
  wire [16:0] _T_379; // @[rvdm.scala 302:30:@315.4]
  wire [29:0] _T_380; // @[rvdm.scala 302:30:@316.4]
  wire [2:0] _T_392; // @[rvdm.scala 309:65:@332.10]
  wire [4:0] abstractcs_datacount; // @[rvdm.scala 498:26:@735.4]
  wire [7:0] _T_398; // @[rvdm.scala 311:46:@345.10]
  wire [2:0] _T_415; // @[rvdm.scala 316:55:@369.8]
  wire  _T_419; // @[rvdm.scala 317:35:@375.8]
  wire  _T_412; // @[rvdm.scala 316:55:@363.8]
  wire  _GEN_5; // @[rvdm.scala 323:44:@389.10]
  wire [1:0] _GEN_12; // @[rvdm.scala 317:44:@376.8]
  wire [2:0] _GEN_0; // @[rvdm.scala 308:36:@324.8]
  wire [2:0] _GEN_2; // @[rvdm.scala 307:43:@323.6]
  wire [2:0] _GEN_20; // @[rvdm.scala 315:40:@355.6]
  wire [2:0] abstractcs_cmderr; // @[rvdm.scala 306:50:@322.4]
  wire [3:0] _T_399; // @[rvdm.scala 311:46:@346.10]
  wire [11:0] _T_400; // @[rvdm.scala 311:46:@347.10]
  wire [11:0] _T_401; // @[rvdm.scala 311:46:@348.10]
  wire [4:0] abstractcs_progbufsize; // @[rvdm.scala 498:26:@735.4]
  wire [7:0] _T_402; // @[rvdm.scala 311:46:@349.10]
  wire [19:0] _T_403; // @[rvdm.scala 311:46:@350.10]
  wire [31:0] _T_404; // @[rvdm.scala 311:46:@351.10]
  wire [31:0] _GEN_1; // @[rvdm.scala 308:36:@324.8]
  wire [31:0] _GEN_3; // @[rvdm.scala 307:43:@323.6]
  wire [15:0] _T_410; // @[rvdm.scala 316:55:@359.8]
  wire  _T_411; // @[rvdm.scala 316:55:@361.8]
  wire  _T_413; // @[rvdm.scala 316:55:@365.8]
  wire  _GEN_9; // @[rvdm.scala 317:44:@376.8]
  wire  _GEN_17; // @[rvdm.scala 315:40:@355.6]
  wire  command_write; // @[rvdm.scala 306:50:@322.4]
  wire [15:0] _GEN_7; // @[rvdm.scala 317:44:@376.8]
  wire [15:0] _GEN_15; // @[rvdm.scala 315:40:@355.6]
  wire [15:0] command_regno; // @[rvdm.scala 306:50:@322.4]
  wire [16:0] _T_420; // @[rvdm.scala 322:40:@381.10]
  wire  _GEN_6; // @[rvdm.scala 317:44:@376.8]
  wire  _GEN_14; // @[rvdm.scala 315:40:@355.6]
  wire  command_postexec; // @[rvdm.scala 306:50:@322.4]
  wire  _GEN_8; // @[rvdm.scala 317:44:@376.8]
  wire  _GEN_16; // @[rvdm.scala 315:40:@355.6]
  wire  command_transfer; // @[rvdm.scala 306:50:@322.4]
  wire [1:0] _T_421; // @[rvdm.scala 322:40:@382.10]
  wire [18:0] _T_422; // @[rvdm.scala 322:40:@383.10]
  wire [3:0] _T_423; // @[rvdm.scala 322:40:@384.10]
  wire [8:0] _T_424; // @[rvdm.scala 322:40:@385.10]
  wire [12:0] _T_425; // @[rvdm.scala 322:40:@386.10]
  wire [31:0] _T_426; // @[rvdm.scala 322:40:@387.10]
  wire [31:0] _GEN_10; // @[rvdm.scala 317:44:@376.8]
  wire  _GEN_11; // @[rvdm.scala 317:44:@376.8]
  wire [31:0] _GEN_13; // @[rvdm.scala 317:44:@376.8]
  wire [31:0] _GEN_18; // @[rvdm.scala 315:40:@355.6]
  wire  _GEN_19; // @[rvdm.scala 315:40:@355.6]
  wire [31:0] _GEN_21; // @[rvdm.scala 315:40:@355.6]
  wire  _T_452; // @[rvdm.scala 342:59:@423.8]
  wire  _T_453; // @[rvdm.scala 342:59:@425.8]
  wire  _T_459; // @[rvdm.scala 342:59:@437.8]
  wire  _GEN_25; // @[rvdm.scala 341:42:@419.6]
  wire  dmcontrol_ndmreset; // @[rvdm.scala 306:50:@322.4]
  wire  _GEN_26; // @[rvdm.scala 341:42:@419.6]
  wire  dmcontrol_dmactive; // @[rvdm.scala 306:50:@322.4]
  wire [1:0] _T_462; // @[rvdm.scala 348:40:@448.8]
  wire [10:0] _T_463; // @[rvdm.scala 348:40:@449.8]
  wire [24:0] _T_464; // @[rvdm.scala 348:40:@450.8]
  wire [26:0] _T_465; // @[rvdm.scala 348:40:@451.8]
  wire [1:0] _T_466; // @[rvdm.scala 348:40:@452.8]
  wire [1:0] _T_467; // @[rvdm.scala 348:40:@453.8]
  wire  _GEN_24; // @[rvdm.scala 341:42:@419.6]
  wire  dmcontrol_hartreset; // @[rvdm.scala 306:50:@322.4]
  wire [2:0] _T_468; // @[rvdm.scala 348:40:@454.8]
  wire [4:0] _T_469; // @[rvdm.scala 348:40:@455.8]
  wire [31:0] _T_470; // @[rvdm.scala 348:40:@456.8]
  wire [31:0] _GEN_27; // @[rvdm.scala 341:42:@419.6]
  wire [2:0] _T_482; // @[rvdm.scala 352:49:@475.8]
  wire  _T_483; // @[rvdm.scala 352:49:@477.8]
  wire [2:0] _T_485; // @[rvdm.scala 352:49:@481.8]
  wire  _T_486; // @[rvdm.scala 352:49:@483.8]
  wire  sbcs_sbaccess32; // @[rvdm.scala 498:26:@735.4]
  wire [1:0] _T_488; // @[rvdm.scala 358:30:@492.8]
  wire [2:0] _T_489; // @[rvdm.scala 358:30:@493.8]
  wire [6:0] sbcs_sbasize; // @[rvdm.scala 498:26:@735.4]
  wire [7:0] _T_490; // @[rvdm.scala 358:30:@494.8]
  wire [8:0] _T_491; // @[rvdm.scala 358:30:@495.8]
  wire [11:0] _T_492; // @[rvdm.scala 358:30:@496.8]
  wire  _GEN_30; // @[rvdm.scala 351:38:@459.6]
  wire  sbcs_sbautoincrement; // @[rvdm.scala 306:50:@322.4]
  wire  _GEN_31; // @[rvdm.scala 351:38:@459.6]
  wire  sbcs_sbautoread; // @[rvdm.scala 306:50:@322.4]
  wire [1:0] _T_493; // @[rvdm.scala 358:30:@497.8]
  wire [2:0] _GEN_32; // @[rvdm.scala 351:38:@459.6]
  wire [2:0] sbcs_sberror; // @[rvdm.scala 306:50:@322.4]
  wire [4:0] _T_494; // @[rvdm.scala 358:30:@498.8]
  wire  _GEN_28; // @[rvdm.scala 351:38:@459.6]
  wire  sbcs_sbsingleread; // @[rvdm.scala 306:50:@322.4]
  wire [11:0] _T_495; // @[rvdm.scala 358:30:@499.8]
  wire [2:0] _GEN_29; // @[rvdm.scala 351:38:@459.6]
  wire [2:0] _GEN_77; // @[rvdm.scala 306:50:@322.4]
  wire [2:0] sbcs_sbaccess; // @[rvdm.scala 498:26:@735.4]
  wire [14:0] _T_496; // @[rvdm.scala 358:30:@500.8]
  wire [19:0] _T_497; // @[rvdm.scala 358:30:@501.8]
  wire [31:0] _T_498; // @[rvdm.scala 358:30:@502.8]
  wire [31:0] _GEN_33; // @[rvdm.scala 351:38:@459.6]
  wire [31:0] _GEN_34; // @[rvdm.scala 362:49:@505.6]
  wire [31:0] _GEN_35; // @[rvdm.scala 362:49:@508.6]
  wire [31:0] _GEN_36; // @[rvdm.scala 362:49:@511.6]
  wire  _GEN_37; // @[rvdm.scala 378:43:@521.8]
  wire  _T_501; // @[rvdm.scala 382:36:@524.8]
  wire [32:0] _T_505; // @[rvdm.scala 387:58:@529.12]
  wire [31:0] _T_506; // @[rvdm.scala 387:58:@530.12]
  wire [31:0] _GEN_38; // @[rvdm.scala 386:44:@528.10]
  wire  _GEN_40; // @[rvdm.scala 382:58:@525.8]
  wire [31:0] _GEN_41; // @[rvdm.scala 382:58:@525.8]
  wire [31:0] _GEN_42; // @[rvdm.scala 368:40:@514.6]
  wire  _GEN_47; // @[rvdm.scala 368:40:@514.6]
  wire  _GEN_48; // @[rvdm.scala 368:40:@514.6]
  wire [31:0] _GEN_49; // @[rvdm.scala 368:40:@514.6]
  wire [31:0] _GEN_50; // @[rvdm.scala 393:44:@535.6]
  wire [31:0] _GEN_51; // @[rvdm.scala 393:44:@538.6]
  wire [31:0] _GEN_52; // @[rvdm.scala 393:44:@541.6]
  wire [31:0] _GEN_53; // @[rvdm.scala 393:44:@544.6]
  wire [31:0] _GEN_54; // @[rvdm.scala 393:44:@547.6]
  wire [31:0] _GEN_55; // @[rvdm.scala 393:44:@550.6]
  wire [31:0] _GEN_56; // @[rvdm.scala 393:44:@553.6]
  wire [31:0] _GEN_57; // @[rvdm.scala 393:44:@556.6]
  wire [31:0] _GEN_58; // @[rvdm.scala 393:44:@559.6]
  wire [31:0] _GEN_59; // @[rvdm.scala 393:44:@562.6]
  wire [31:0] _GEN_60; // @[rvdm.scala 393:44:@565.6]
  wire [31:0] _GEN_61; // @[rvdm.scala 393:44:@568.6]
  wire [31:0] _GEN_63; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_68; // @[rvdm.scala 306:50:@322.4]
  wire  _GEN_69; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_75; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_81; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_82; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_83; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_84; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_85; // @[rvdm.scala 306:50:@322.4]
  wire  _GEN_90; // @[rvdm.scala 306:50:@322.4]
  wire  _GEN_91; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_92; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_93; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_94; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_95; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_96; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_97; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_98; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_99; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_100; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_101; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_102; // @[rvdm.scala 306:50:@322.4]
  wire [31:0] _GEN_103; // @[rvdm.scala 306:50:@322.4]
  wire  _T_514; // @[Mux.scala 46:19:@578.4]
  wire [31:0] _T_515; // @[Mux.scala 46:16:@579.4]
  wire  _T_516; // @[Mux.scala 46:19:@580.4]
  wire [31:0] _T_517; // @[Mux.scala 46:16:@581.4]
  wire  _T_518; // @[Mux.scala 46:19:@582.4]
  wire [31:0] _T_519; // @[Mux.scala 46:16:@583.4]
  wire  _T_520; // @[Mux.scala 46:19:@584.4]
  wire [31:0] _T_521; // @[Mux.scala 46:16:@585.4]
  wire  _T_522; // @[Mux.scala 46:19:@586.4]
  wire [31:0] _T_523; // @[Mux.scala 46:16:@587.4]
  wire  _T_524; // @[Mux.scala 46:19:@588.4]
  wire [31:0] _T_525; // @[Mux.scala 46:16:@589.4]
  wire  _T_526; // @[Mux.scala 46:19:@590.4]
  wire [31:0] _T_527; // @[Mux.scala 46:16:@591.4]
  wire  _T_528; // @[Mux.scala 46:19:@592.4]
  wire [31:0] _T_529; // @[Mux.scala 46:16:@593.4]
  wire  _T_530; // @[Mux.scala 46:19:@594.4]
  wire [31:0] _T_531; // @[Mux.scala 46:16:@595.4]
  wire  _T_532; // @[Mux.scala 46:19:@596.4]
  wire [31:0] _T_533; // @[Mux.scala 46:16:@597.4]
  wire  _T_534; // @[Mux.scala 46:19:@598.4]
  wire [31:0] _T_535; // @[Mux.scala 46:16:@599.4]
  wire  _T_536; // @[Mux.scala 46:19:@600.4]
  wire [31:0] _T_537; // @[Mux.scala 46:16:@601.4]
  wire  _T_538; // @[Mux.scala 46:19:@602.4]
  wire [31:0] _T_539; // @[Mux.scala 46:16:@603.4]
  wire  _T_540; // @[Mux.scala 46:19:@604.4]
  wire [31:0] _T_541; // @[Mux.scala 46:16:@605.4]
  wire  _T_542; // @[Mux.scala 46:19:@606.4]
  wire [31:0] _T_543; // @[Mux.scala 46:16:@607.4]
  wire  _T_544; // @[Mux.scala 46:19:@608.4]
  wire [31:0] _T_545; // @[Mux.scala 46:16:@609.4]
  wire  _T_546; // @[Mux.scala 46:19:@610.4]
  wire [31:0] _T_547; // @[Mux.scala 46:16:@611.4]
  wire  _T_548; // @[Mux.scala 46:19:@612.4]
  wire [31:0] _T_549; // @[Mux.scala 46:16:@613.4]
  wire  _T_550; // @[Mux.scala 46:19:@614.4]
  wire [31:0] _T_551; // @[Mux.scala 46:16:@615.4]
  wire  _T_552; // @[Mux.scala 46:19:@616.4]
  wire [31:0] _T_553; // @[Mux.scala 46:16:@617.4]
  wire  _T_554; // @[Mux.scala 46:19:@618.4]
  wire [31:0] _T_555; // @[Mux.scala 46:16:@619.4]
  wire  _T_556; // @[Mux.scala 46:19:@620.4]
  wire [31:0] _T_557; // @[Mux.scala 46:16:@621.4]
  wire  _T_558; // @[Mux.scala 46:19:@622.4]
  wire [31:0] _T_559; // @[Mux.scala 46:16:@623.4]
  wire  _T_560; // @[Mux.scala 46:19:@624.4]
  wire [31:0] _T_561; // @[Mux.scala 46:16:@625.4]
  wire  _T_562; // @[Mux.scala 46:19:@626.4]
  wire [31:0] _T_563; // @[Mux.scala 46:16:@627.4]
  wire  _T_564; // @[Mux.scala 46:19:@628.4]
  wire [31:0] _T_565; // @[Mux.scala 46:16:@629.4]
  wire  _T_566; // @[Mux.scala 46:19:@630.4]
  wire [31:0] _T_567; // @[Mux.scala 46:16:@631.4]
  wire  _T_568; // @[Mux.scala 46:19:@632.4]
  wire [31:0] _T_569; // @[Mux.scala 46:16:@633.4]
  wire  _T_570; // @[Mux.scala 46:19:@634.4]
  wire [31:0] _T_571; // @[Mux.scala 46:16:@635.4]
  wire  _T_572; // @[Mux.scala 46:19:@636.4]
  wire [31:0] _T_573; // @[Mux.scala 46:16:@637.4]
  wire  _T_574; // @[Mux.scala 46:19:@638.4]
  wire [31:0] _T_575; // @[Mux.scala 46:16:@639.4]
  wire  _T_576; // @[Mux.scala 46:19:@640.4]
  wire [31:0] _T_577; // @[Mux.scala 46:16:@641.4]
  wire  _T_578; // @[Mux.scala 46:19:@642.4]
  wire [31:0] _T_579; // @[Mux.scala 46:16:@643.4]
  wire  _T_580; // @[Mux.scala 46:19:@644.4]
  wire [31:0] _T_581; // @[Mux.scala 46:16:@645.4]
  wire  _T_582; // @[Mux.scala 46:19:@646.4]
  wire [31:0] _T_583; // @[Mux.scala 46:16:@647.4]
  wire  _T_584; // @[Mux.scala 46:19:@648.4]
  wire [31:0] _T_585; // @[Mux.scala 46:16:@649.4]
  wire  _T_586; // @[Mux.scala 46:19:@650.4]
  wire [31:0] _T_587; // @[Mux.scala 46:16:@651.4]
  wire  _T_588; // @[Mux.scala 46:19:@652.4]
  wire [31:0] _T_589; // @[Mux.scala 46:16:@653.4]
  wire  _T_590; // @[Mux.scala 46:19:@654.4]
  wire [31:0] _T_591; // @[Mux.scala 46:16:@655.4]
  wire  _T_592; // @[Mux.scala 46:19:@656.4]
  wire [31:0] _T_593; // @[Mux.scala 46:16:@657.4]
  wire  _T_594; // @[Mux.scala 46:19:@658.4]
  wire [31:0] _T_595; // @[Mux.scala 46:16:@659.4]
  wire  _T_596; // @[Mux.scala 46:19:@660.4]
  wire [31:0] _T_597; // @[Mux.scala 46:16:@661.4]
  wire  _T_598; // @[Mux.scala 46:19:@662.4]
  wire [31:0] _T_599; // @[Mux.scala 46:16:@663.4]
  wire  _T_600; // @[Mux.scala 46:19:@664.4]
  wire [31:0] _T_601; // @[Mux.scala 46:16:@665.4]
  wire [15:0] _T_604; // @[rvdm.scala 404:38:@668.4]
  wire [4:0] _T_605; // @[rvdm.scala 404:47:@669.4]
  wire  cmd_regrw; // @[rvdm.scala 406:39:@671.4]
  wire [31:0] _GEN_106; // @[rvdm.scala 408:29:@673.6]
  wire  _GEN_108; // @[rvdm.scala 407:21:@672.4]
  wire [31:0] _GEN_109; // @[rvdm.scala 407:21:@672.4]
  wire  _GEN_110; // @[rvdm.scala 407:21:@672.4]
  wire  _T_608; // @[rvdm.scala 424:29:@682.4]
  wire  _T_609; // @[rvdm.scala 424:47:@683.4]
  wire  _T_611; // @[rvdm.scala 434:37:@690.8]
  wire [31:0] _GEN_111; // @[rvdm.scala 441:44:@696.10]
  wire [31:0] _GEN_113; // @[rvdm.scala 434:59:@691.8]
  wire  _GEN_114; // @[rvdm.scala 434:59:@691.8]
  wire  _GEN_115; // @[rvdm.scala 434:59:@691.8]
  wire  _GEN_116; // @[rvdm.scala 434:59:@691.8]
  wire [31:0] _GEN_117; // @[rvdm.scala 434:59:@691.8]
  wire  _GEN_118; // @[rvdm.scala 455:38:@711.8]
  wire  _GEN_119; // @[rvdm.scala 432:36:@688.6]
  wire [31:0] _GEN_120; // @[rvdm.scala 432:36:@688.6]
  wire  _GEN_121; // @[rvdm.scala 432:36:@688.6]
  wire  _GEN_122; // @[rvdm.scala 432:36:@688.6]
  wire [31:0] _GEN_123; // @[rvdm.scala 432:36:@688.6]
  wire  _GEN_124; // @[rvdm.scala 424:74:@684.4]
  wire  _GEN_127; // @[rvdm.scala 424:74:@684.4]
  wire [31:0] _GEN_128; // @[rvdm.scala 424:74:@684.4]
  wire  _GEN_129; // @[rvdm.scala 424:74:@684.4]
  wire  _GEN_130; // @[rvdm.scala 424:74:@684.4]
  wire [31:0] _GEN_131; // @[rvdm.scala 424:74:@684.4]
  wire  _T_623; // @[rvdm.scala 463:10:@716.4]
  wire  _GEN_132; // @[rvdm.scala 463:39:@717.4]
  wire  _T_625; // @[rvdm.scala 479:29:@720.4]
  wire  _T_627; // @[rvdm.scala 490:32:@724.4]
  wire  _T_628; // @[rvdm.scala 490:45:@725.4]
  wire  _GEN_133; // @[rvdm.scala 490:65:@726.4]
  wire  _T_631; // @[rvdm.scala 493:32:@729.4]
  wire  _T_632; // @[rvdm.scala 493:45:@730.4]
  wire  _GEN_134; // @[rvdm.scala 493:65:@731.4]
  wire [31:0] _GEN_135; // @[rvdm.scala 498:26:@735.4]
  wire [31:0] _GEN_136; // @[rvdm.scala 498:26:@735.4]
  wire [31:0] _GEN_137; // @[rvdm.scala 498:26:@735.4]
  wire [31:0] _GEN_138; // @[rvdm.scala 498:26:@735.4]
  wire [31:0] _GEN_139; // @[rvdm.scala 498:26:@735.4]
  wire [31:0] _GEN_140; // @[rvdm.scala 498:26:@735.4]
  wire [31:0] _GEN_141; // @[rvdm.scala 498:26:@735.4]
  wire  _GEN_142; // @[rvdm.scala 498:26:@735.4]
  wire  _GEN_143; // @[rvdm.scala 498:26:@735.4]
  wire [29:0] _GEN_146; // @[rvdm.scala 498:26:@735.4]
  wire [31:0] _GEN_152; // @[rvdm.scala 498:26:@735.4]
  wire  _GEN_153; // @[rvdm.scala 498:26:@735.4]
  wire  _GEN_154; // @[rvdm.scala 498:26:@735.4]
  wire [1:0] _GEN_155; // @[rvdm.scala 498:26:@735.4]
  wire  _GEN_156; // @[rvdm.scala 498:26:@735.4]
  wire  _GEN_157; // @[rvdm.scala 498:26:@735.4]
  assign _T_132 = io_dmi_req_bits_addr == 7'h10; // @[rvdm.scala 278:74:@51.4]
  assign _T_144 = io_dmi_req_bits_addr == 7'h16; // @[rvdm.scala 278:74:@57.4]
  assign _T_146 = io_dmi_req_bits_addr == 7'h17; // @[rvdm.scala 278:74:@58.4]
  assign _T_154 = io_dmi_req_bits_addr == 7'h38; // @[rvdm.scala 278:74:@62.4]
  assign _T_156 = io_dmi_req_bits_addr == 7'h4; // @[rvdm.scala 278:74:@63.4]
  assign _T_158 = io_dmi_req_bits_addr == 7'h5; // @[rvdm.scala 278:74:@64.4]
  assign _T_160 = io_dmi_req_bits_addr == 7'h6; // @[rvdm.scala 278:74:@65.4]
  assign _T_162 = io_dmi_req_bits_addr == 7'h7; // @[rvdm.scala 278:74:@66.4]
  assign _T_164 = io_dmi_req_bits_addr == 7'h8; // @[rvdm.scala 278:74:@67.4]
  assign _T_166 = io_dmi_req_bits_addr == 7'h9; // @[rvdm.scala 278:74:@68.4]
  assign _T_168 = io_dmi_req_bits_addr == 7'ha; // @[rvdm.scala 278:74:@69.4]
  assign _T_170 = io_dmi_req_bits_addr == 7'hb; // @[rvdm.scala 278:74:@70.4]
  assign _T_172 = io_dmi_req_bits_addr == 7'hc; // @[rvdm.scala 278:74:@71.4]
  assign _T_174 = io_dmi_req_bits_addr == 7'hd; // @[rvdm.scala 278:74:@72.4]
  assign _T_176 = io_dmi_req_bits_addr == 7'he; // @[rvdm.scala 278:74:@73.4]
  assign _T_178 = io_dmi_req_bits_addr == 7'hf; // @[rvdm.scala 278:74:@74.4]
  assign _T_212 = io_dmi_req_bits_addr == 7'h39; // @[rvdm.scala 278:74:@91.4]
  assign _T_214 = io_dmi_req_bits_addr == 7'h3a; // @[rvdm.scala 278:74:@92.4]
  assign _T_216 = io_dmi_req_bits_addr == 7'h3b; // @[rvdm.scala 278:74:@93.4]
  assign _T_218 = io_dmi_req_bits_addr == 7'h3c; // @[rvdm.scala 278:74:@94.4]
  assign _T_277 = reg_dmstatus[29:0]; // @[:@100.4]
  assign _T_278 = _T_277[3:0]; // @[rvdm.scala 290:42:@102.4]
  assign dmstatus_devtreevalid = _T_277[4]; // @[rvdm.scala 290:42:@104.4]
  assign dmstatus_rsrvd4 = _T_277[5]; // @[rvdm.scala 290:42:@106.4]
  assign dmstatus_authbusy = _T_277[6]; // @[rvdm.scala 290:42:@108.4]
  assign _T_282 = _T_277[7]; // @[rvdm.scala 290:42:@110.4]
  assign dmstatus_anyhalted = _T_277[8]; // @[rvdm.scala 290:42:@112.4]
  assign dmstatus_anyrunning = _T_277[10]; // @[rvdm.scala 290:42:@116.4]
  assign dmstatus_anyunavail = _T_277[12]; // @[rvdm.scala 290:42:@120.4]
  assign dmstatus_allunavail = _T_277[13]; // @[rvdm.scala 290:42:@122.4]
  assign dmstatus_anynonexistent = _T_277[14]; // @[rvdm.scala 290:42:@124.4]
  assign dmstatus_allnonexistent = _T_277[15]; // @[rvdm.scala 290:42:@126.4]
  assign dmstatus_allresumeack = _T_277[16]; // @[rvdm.scala 290:42:@128.4]
  assign dmstatus_anyhavereset = _T_277[17]; // @[rvdm.scala 290:42:@130.4]
  assign dmstatus_allhavereset = _T_277[18]; // @[rvdm.scala 290:42:@132.4]
  assign dmstatus_rsrvd3 = _T_277[19]; // @[rvdm.scala 290:42:@134.4]
  assign dmstatus_impebreak = _T_277[20]; // @[rvdm.scala 290:42:@136.4]
  assign dmstatus_rsrvd2 = _T_277[21]; // @[rvdm.scala 290:42:@138.4]
  assign dmstatus_dmerr = _T_277[24:22]; // @[rvdm.scala 290:42:@140.4]
  assign dmstatus_rsrvd1 = _T_277[29:25]; // @[rvdm.scala 290:42:@142.4]
  assign _T_305 = reg_dmcontrol[0]; // @[rvdm.scala 292:44:@169.4]
  assign _T_306 = reg_dmcontrol[1]; // @[rvdm.scala 292:44:@171.4]
  assign dmcontrol_rsrvd2 = reg_dmcontrol[15:2]; // @[rvdm.scala 292:44:@173.4]
  assign dmcontrol_hartsel = reg_dmcontrol[25:16]; // @[rvdm.scala 292:44:@175.4]
  assign dmcontrol_hasel = reg_dmcontrol[26]; // @[rvdm.scala 292:44:@177.4]
  assign dmcontrol_rsrvd1 = reg_dmcontrol[27]; // @[rvdm.scala 292:44:@179.4]
  assign dmcontrol_ackharvereset = reg_dmcontrol[28]; // @[rvdm.scala 292:44:@181.4]
  assign _T_312 = reg_dmcontrol[29]; // @[rvdm.scala 292:44:@183.4]
  assign _T_313 = reg_dmcontrol[30]; // @[rvdm.scala 292:44:@185.4]
  assign _T_314 = reg_dmcontrol[31]; // @[rvdm.scala 292:44:@187.4]
  assign sbcs_sbaccess8 = reg_sbcs[0]; // @[rvdm.scala 294:34:@203.4]
  assign sbcs_sbaccess16 = reg_sbcs[1]; // @[rvdm.scala 294:34:@205.4]
  assign _T_323 = reg_sbcs[2]; // @[rvdm.scala 294:34:@207.4]
  assign sbcs_sbaccess64 = reg_sbcs[3]; // @[rvdm.scala 294:34:@209.4]
  assign sbcs_sbaccess128 = reg_sbcs[4]; // @[rvdm.scala 294:34:@211.4]
  assign _T_326 = reg_sbcs[11:5]; // @[rvdm.scala 294:34:@213.4]
  assign _T_327 = reg_sbcs[14:12]; // @[rvdm.scala 294:34:@215.4]
  assign _T_328 = reg_sbcs[15]; // @[rvdm.scala 294:34:@217.4]
  assign _T_329 = reg_sbcs[16]; // @[rvdm.scala 294:34:@219.4]
  assign _T_330 = reg_sbcs[19:17]; // @[rvdm.scala 294:34:@221.4]
  assign _T_331 = reg_sbcs[20]; // @[rvdm.scala 294:34:@223.4]
  assign sbcs_rsrvd1 = reg_sbcs[31:21]; // @[rvdm.scala 294:34:@225.4]
  assign _T_339 = reg_abstractcs[4:0]; // @[rvdm.scala 296:46:@243.4]
  assign abstractcs_rsrvd4 = reg_abstractcs[7:5]; // @[rvdm.scala 296:46:@245.4]
  assign _T_341 = reg_abstractcs[10:8]; // @[rvdm.scala 296:46:@247.4]
  assign abstractcs_rsrvd3 = reg_abstractcs[11]; // @[rvdm.scala 296:46:@249.4]
  assign abstractcs_busy = reg_abstractcs[12]; // @[rvdm.scala 296:46:@251.4]
  assign abstractcs_rsrvd2 = reg_abstractcs[23:13]; // @[rvdm.scala 296:46:@253.4]
  assign _T_345 = reg_abstractcs[28:24]; // @[rvdm.scala 296:46:@255.4]
  assign abstractcs_rsrvd1 = reg_abstractcs[31:29]; // @[rvdm.scala 296:46:@257.4]
  assign _T_353 = reg_command[15:0]; // @[rvdm.scala 298:40:@271.4]
  assign _T_354 = reg_command[16]; // @[rvdm.scala 298:40:@273.4]
  assign _T_355 = reg_command[17]; // @[rvdm.scala 298:40:@275.4]
  assign _T_356 = reg_command[18]; // @[rvdm.scala 298:40:@277.4]
  assign command_rsrvd2 = reg_command[19]; // @[rvdm.scala 298:40:@279.4]
  assign command_size = reg_command[22:20]; // @[rvdm.scala 298:40:@281.4]
  assign command_rsrvd1 = reg_command[23]; // @[rvdm.scala 298:40:@283.4]
  assign command_cmdtype = reg_command[31:24]; // @[rvdm.scala 298:40:@285.4]
  assign dmstatus_version = reset ? 4'h2 : _T_278; // @[rvdm.scala 498:26:@735.4]
  assign _T_361 = {dmstatus_devtreevalid,dmstatus_version}; // @[rvdm.scala 302:30:@297.4]
  assign dmstatus_authenticated = reset ? 1'h1 : _T_282; // @[rvdm.scala 498:26:@735.4]
  assign _T_362 = {dmstatus_authenticated,dmstatus_authbusy}; // @[rvdm.scala 302:30:@298.4]
  assign _T_363 = {_T_362,dmstatus_rsrvd4}; // @[rvdm.scala 302:30:@299.4]
  assign _T_364 = {_T_363,_T_361}; // @[rvdm.scala 302:30:@300.4]
  assign _T_384 = io_dmi_req_bits_op == 2'h2; // @[rvdm.scala 306:29:@321.4]
  assign _T_461 = io_dmi_req_bits_data[31]; // @[rvdm.scala 342:59:@441.8]
  assign _GEN_22 = _T_132 ? _T_461 : _T_314; // @[rvdm.scala 341:42:@419.6]
  assign dmcontrol_haltreq = _T_384 ? _GEN_22 : _T_314; // @[rvdm.scala 306:50:@322.4]
  assign _T_365 = {dmcontrol_haltreq,dmstatus_anyhalted}; // @[rvdm.scala 302:30:@301.4]
  assign _T_460 = io_dmi_req_bits_data[30]; // @[rvdm.scala 342:59:@439.8]
  assign _GEN_23 = _T_132 ? _T_460 : _T_313; // @[rvdm.scala 341:42:@419.6]
  assign dmcontrol_resumereq = _T_384 ? _GEN_23 : _T_313; // @[rvdm.scala 306:50:@322.4]
  assign _T_366 = {dmstatus_anyunavail,dmcontrol_resumereq}; // @[rvdm.scala 302:30:@302.4]
  assign _T_367 = {_T_366,dmstatus_anyrunning}; // @[rvdm.scala 302:30:@303.4]
  assign _T_368 = {_T_367,_T_365}; // @[rvdm.scala 302:30:@304.4]
  assign _T_369 = {_T_368,_T_364}; // @[rvdm.scala 302:30:@305.4]
  assign _T_370 = {dmstatus_anynonexistent,dmstatus_allunavail}; // @[rvdm.scala 302:30:@306.4]
  assign _T_371 = {dmstatus_anyhavereset,dmstatus_allresumeack}; // @[rvdm.scala 302:30:@307.4]
  assign _T_372 = {_T_371,dmstatus_allnonexistent}; // @[rvdm.scala 302:30:@308.4]
  assign _T_373 = {_T_372,_T_370}; // @[rvdm.scala 302:30:@309.4]
  assign _T_374 = {dmstatus_impebreak,dmstatus_rsrvd3}; // @[rvdm.scala 302:30:@310.4]
  assign _T_375 = {_T_374,dmstatus_allhavereset}; // @[rvdm.scala 302:30:@311.4]
  assign _T_376 = {dmstatus_rsrvd1,dmstatus_dmerr}; // @[rvdm.scala 302:30:@312.4]
  assign _T_377 = {_T_376,dmstatus_rsrvd2}; // @[rvdm.scala 302:30:@313.4]
  assign _T_378 = {_T_377,_T_375}; // @[rvdm.scala 302:30:@314.4]
  assign _T_379 = {_T_378,_T_373}; // @[rvdm.scala 302:30:@315.4]
  assign _T_380 = {_T_379,_T_369}; // @[rvdm.scala 302:30:@316.4]
  assign _T_392 = io_dmi_req_bits_data[10:8]; // @[rvdm.scala 309:65:@332.10]
  assign abstractcs_datacount = reset ? 5'hc : _T_339; // @[rvdm.scala 498:26:@735.4]
  assign _T_398 = {abstractcs_rsrvd4,abstractcs_datacount}; // @[rvdm.scala 311:46:@345.10]
  assign _T_415 = io_dmi_req_bits_data[22:20]; // @[rvdm.scala 316:55:@369.8]
  assign _T_419 = _T_415 == 3'h2; // @[rvdm.scala 317:35:@375.8]
  assign _T_412 = io_dmi_req_bits_data[17]; // @[rvdm.scala 316:55:@363.8]
  assign _GEN_5 = _T_412 ? 1'h0 : 1'h1; // @[rvdm.scala 323:44:@389.10]
  assign _GEN_12 = _T_419 ? {{1'd0}, _GEN_5} : 2'h2; // @[rvdm.scala 317:44:@376.8]
  assign _GEN_0 = io_dmi_req_valid ? _T_392 : _T_341; // @[rvdm.scala 308:36:@324.8]
  assign _GEN_2 = _T_144 ? _GEN_0 : _T_341; // @[rvdm.scala 307:43:@323.6]
  assign _GEN_20 = _T_146 ? {{1'd0}, _GEN_12} : _GEN_2; // @[rvdm.scala 315:40:@355.6]
  assign abstractcs_cmderr = _T_384 ? _GEN_20 : _T_341; // @[rvdm.scala 306:50:@322.4]
  assign _T_399 = {abstractcs_rsrvd3,abstractcs_cmderr}; // @[rvdm.scala 311:46:@346.10]
  assign _T_400 = {_T_399,_T_398}; // @[rvdm.scala 311:46:@347.10]
  assign _T_401 = {abstractcs_rsrvd2,abstractcs_busy}; // @[rvdm.scala 311:46:@348.10]
  assign abstractcs_progbufsize = reset ? 5'h10 : _T_345; // @[rvdm.scala 498:26:@735.4]
  assign _T_402 = {abstractcs_rsrvd1,abstractcs_progbufsize}; // @[rvdm.scala 311:46:@349.10]
  assign _T_403 = {_T_402,_T_401}; // @[rvdm.scala 311:46:@350.10]
  assign _T_404 = {_T_403,_T_400}; // @[rvdm.scala 311:46:@351.10]
  assign _GEN_1 = io_dmi_req_valid ? _T_404 : reg_abstractcs; // @[rvdm.scala 308:36:@324.8]
  assign _GEN_3 = _T_144 ? _GEN_1 : reg_abstractcs; // @[rvdm.scala 307:43:@323.6]
  assign _T_410 = io_dmi_req_bits_data[15:0]; // @[rvdm.scala 316:55:@359.8]
  assign _T_411 = io_dmi_req_bits_data[16]; // @[rvdm.scala 316:55:@361.8]
  assign _T_413 = io_dmi_req_bits_data[18]; // @[rvdm.scala 316:55:@365.8]
  assign _GEN_9 = _T_419 ? _T_411 : _T_354; // @[rvdm.scala 317:44:@376.8]
  assign _GEN_17 = _T_146 ? _GEN_9 : _T_354; // @[rvdm.scala 315:40:@355.6]
  assign command_write = _T_384 ? _GEN_17 : _T_354; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_7 = _T_419 ? _T_410 : _T_353; // @[rvdm.scala 317:44:@376.8]
  assign _GEN_15 = _T_146 ? _GEN_7 : _T_353; // @[rvdm.scala 315:40:@355.6]
  assign command_regno = _T_384 ? _GEN_15 : _T_353; // @[rvdm.scala 306:50:@322.4]
  assign _T_420 = {command_write,command_regno}; // @[rvdm.scala 322:40:@381.10]
  assign _GEN_6 = _T_419 ? _T_413 : _T_356; // @[rvdm.scala 317:44:@376.8]
  assign _GEN_14 = _T_146 ? _GEN_6 : _T_356; // @[rvdm.scala 315:40:@355.6]
  assign command_postexec = _T_384 ? _GEN_14 : _T_356; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_8 = _T_419 ? _T_412 : _T_355; // @[rvdm.scala 317:44:@376.8]
  assign _GEN_16 = _T_146 ? _GEN_8 : _T_355; // @[rvdm.scala 315:40:@355.6]
  assign command_transfer = _T_384 ? _GEN_16 : _T_355; // @[rvdm.scala 306:50:@322.4]
  assign _T_421 = {command_postexec,command_transfer}; // @[rvdm.scala 322:40:@382.10]
  assign _T_422 = {_T_421,_T_420}; // @[rvdm.scala 322:40:@383.10]
  assign _T_423 = {command_size,command_rsrvd2}; // @[rvdm.scala 322:40:@384.10]
  assign _T_424 = {command_cmdtype,command_rsrvd1}; // @[rvdm.scala 322:40:@385.10]
  assign _T_425 = {_T_424,_T_423}; // @[rvdm.scala 322:40:@386.10]
  assign _T_426 = {_T_425,_T_422}; // @[rvdm.scala 322:40:@387.10]
  assign _GEN_10 = _T_419 ? _T_426 : reg_command; // @[rvdm.scala 317:44:@376.8]
  assign _GEN_11 = _T_419 ? _T_412 : 1'h0; // @[rvdm.scala 317:44:@376.8]
  assign _GEN_13 = _T_419 ? _T_404 : _T_404; // @[rvdm.scala 317:44:@376.8]
  assign _GEN_18 = _T_146 ? _GEN_10 : reg_command; // @[rvdm.scala 315:40:@355.6]
  assign _GEN_19 = _T_146 ? _GEN_11 : reg_regrw; // @[rvdm.scala 315:40:@355.6]
  assign _GEN_21 = _T_146 ? _GEN_13 : _GEN_3; // @[rvdm.scala 315:40:@355.6]
  assign _T_452 = io_dmi_req_bits_data[0]; // @[rvdm.scala 342:59:@423.8]
  assign _T_453 = io_dmi_req_bits_data[1]; // @[rvdm.scala 342:59:@425.8]
  assign _T_459 = io_dmi_req_bits_data[29]; // @[rvdm.scala 342:59:@437.8]
  assign _GEN_25 = _T_132 ? _T_453 : _T_306; // @[rvdm.scala 341:42:@419.6]
  assign dmcontrol_ndmreset = _T_384 ? _GEN_25 : _T_306; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_26 = _T_132 ? _T_452 : _T_305; // @[rvdm.scala 341:42:@419.6]
  assign dmcontrol_dmactive = _T_384 ? _GEN_26 : _T_305; // @[rvdm.scala 306:50:@322.4]
  assign _T_462 = {dmcontrol_ndmreset,dmcontrol_dmactive}; // @[rvdm.scala 348:40:@448.8]
  assign _T_463 = {dmcontrol_hasel,dmcontrol_hartsel}; // @[rvdm.scala 348:40:@449.8]
  assign _T_464 = {_T_463,dmcontrol_rsrvd2}; // @[rvdm.scala 348:40:@450.8]
  assign _T_465 = {_T_464,_T_462}; // @[rvdm.scala 348:40:@451.8]
  assign _T_466 = {dmcontrol_ackharvereset,dmcontrol_rsrvd1}; // @[rvdm.scala 348:40:@452.8]
  assign _T_467 = {dmcontrol_haltreq,dmcontrol_resumereq}; // @[rvdm.scala 348:40:@453.8]
  assign _GEN_24 = _T_132 ? _T_459 : _T_312; // @[rvdm.scala 341:42:@419.6]
  assign dmcontrol_hartreset = _T_384 ? _GEN_24 : _T_312; // @[rvdm.scala 306:50:@322.4]
  assign _T_468 = {_T_467,dmcontrol_hartreset}; // @[rvdm.scala 348:40:@454.8]
  assign _T_469 = {_T_468,_T_466}; // @[rvdm.scala 348:40:@455.8]
  assign _T_470 = {_T_469,_T_465}; // @[rvdm.scala 348:40:@456.8]
  assign _GEN_27 = _T_132 ? _T_470 : reg_dmcontrol; // @[rvdm.scala 341:42:@419.6]
  assign _T_482 = io_dmi_req_bits_data[14:12]; // @[rvdm.scala 352:49:@475.8]
  assign _T_483 = io_dmi_req_bits_data[15]; // @[rvdm.scala 352:49:@477.8]
  assign _T_485 = io_dmi_req_bits_data[19:17]; // @[rvdm.scala 352:49:@481.8]
  assign _T_486 = io_dmi_req_bits_data[20]; // @[rvdm.scala 352:49:@483.8]
  assign sbcs_sbaccess32 = reset ? 1'h1 : _T_323; // @[rvdm.scala 498:26:@735.4]
  assign _T_488 = {sbcs_sbaccess32,sbcs_sbaccess16}; // @[rvdm.scala 358:30:@492.8]
  assign _T_489 = {_T_488,sbcs_sbaccess8}; // @[rvdm.scala 358:30:@493.8]
  assign sbcs_sbasize = reset ? 7'h20 : _T_326; // @[rvdm.scala 498:26:@735.4]
  assign _T_490 = {sbcs_sbasize,sbcs_sbaccess128}; // @[rvdm.scala 358:30:@494.8]
  assign _T_491 = {_T_490,sbcs_sbaccess64}; // @[rvdm.scala 358:30:@495.8]
  assign _T_492 = {_T_491,_T_489}; // @[rvdm.scala 358:30:@496.8]
  assign _GEN_30 = _T_154 ? _T_411 : _T_329; // @[rvdm.scala 351:38:@459.6]
  assign sbcs_sbautoincrement = _T_384 ? _GEN_30 : _T_329; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_31 = _T_154 ? _T_483 : _T_328; // @[rvdm.scala 351:38:@459.6]
  assign sbcs_sbautoread = _T_384 ? _GEN_31 : _T_328; // @[rvdm.scala 306:50:@322.4]
  assign _T_493 = {sbcs_sbautoincrement,sbcs_sbautoread}; // @[rvdm.scala 358:30:@497.8]
  assign _GEN_32 = _T_154 ? _T_482 : _T_327; // @[rvdm.scala 351:38:@459.6]
  assign sbcs_sberror = _T_384 ? _GEN_32 : _T_327; // @[rvdm.scala 306:50:@322.4]
  assign _T_494 = {_T_493,sbcs_sberror}; // @[rvdm.scala 358:30:@498.8]
  assign _GEN_28 = _T_154 ? _T_486 : _T_331; // @[rvdm.scala 351:38:@459.6]
  assign sbcs_sbsingleread = _T_384 ? _GEN_28 : _T_331; // @[rvdm.scala 306:50:@322.4]
  assign _T_495 = {sbcs_rsrvd1,sbcs_sbsingleread}; // @[rvdm.scala 358:30:@499.8]
  assign _GEN_29 = _T_154 ? _T_485 : _T_330; // @[rvdm.scala 351:38:@459.6]
  assign _GEN_77 = _T_384 ? _GEN_29 : _T_330; // @[rvdm.scala 306:50:@322.4]
  assign sbcs_sbaccess = reset ? 3'h2 : _GEN_77; // @[rvdm.scala 498:26:@735.4]
  assign _T_496 = {_T_495,sbcs_sbaccess}; // @[rvdm.scala 358:30:@500.8]
  assign _T_497 = {_T_496,_T_494}; // @[rvdm.scala 358:30:@501.8]
  assign _T_498 = {_T_497,_T_492}; // @[rvdm.scala 358:30:@502.8]
  assign _GEN_33 = _T_154 ? _T_498 : reg_sbcs; // @[rvdm.scala 351:38:@459.6]
  assign _GEN_34 = _T_212 ? io_dmi_req_bits_data : reg_sbaddress_0; // @[rvdm.scala 362:49:@505.6]
  assign _GEN_35 = _T_214 ? io_dmi_req_bits_data : reg_sbaddress_1; // @[rvdm.scala 362:49:@508.6]
  assign _GEN_36 = _T_216 ? io_dmi_req_bits_data : reg_sbaddress_2; // @[rvdm.scala 362:49:@511.6]
  assign _GEN_37 = reg_delay_mrwdata_valid ? 1'h0 : 1'h1; // @[rvdm.scala 378:43:@521.8]
  assign _T_501 = io_ddmem_req_ready & reg_ddmem_req_valid; // @[rvdm.scala 382:36:@524.8]
  assign _T_505 = reg_sbaddress_0 + 32'h4; // @[rvdm.scala 387:58:@529.12]
  assign _T_506 = _T_505[31:0]; // @[rvdm.scala 387:58:@530.12]
  assign _GEN_38 = sbcs_sbautoincrement ? _T_506 : _GEN_34; // @[rvdm.scala 386:44:@528.10]
  assign _GEN_40 = _T_501 ? 1'h0 : _GEN_37; // @[rvdm.scala 382:58:@525.8]
  assign _GEN_41 = _T_501 ? _GEN_38 : _GEN_34; // @[rvdm.scala 382:58:@525.8]
  assign _GEN_42 = _T_218 ? io_dmi_req_bits_data : reg_sbdata_0; // @[rvdm.scala 368:40:@514.6]
  assign _GEN_47 = _T_218 ? _GEN_40 : 1'h0; // @[rvdm.scala 368:40:@514.6]
  assign _GEN_48 = _T_218 ? _T_501 : 1'h0; // @[rvdm.scala 368:40:@514.6]
  assign _GEN_49 = _T_218 ? _GEN_41 : _GEN_34; // @[rvdm.scala 368:40:@514.6]
  assign _GEN_50 = _T_156 ? io_dmi_req_bits_data : reg_data_0; // @[rvdm.scala 393:44:@535.6]
  assign _GEN_51 = _T_158 ? io_dmi_req_bits_data : reg_data_1; // @[rvdm.scala 393:44:@538.6]
  assign _GEN_52 = _T_160 ? io_dmi_req_bits_data : reg_data_2; // @[rvdm.scala 393:44:@541.6]
  assign _GEN_53 = _T_162 ? io_dmi_req_bits_data : reg_data_3; // @[rvdm.scala 393:44:@544.6]
  assign _GEN_54 = _T_164 ? io_dmi_req_bits_data : reg_data_4; // @[rvdm.scala 393:44:@547.6]
  assign _GEN_55 = _T_166 ? io_dmi_req_bits_data : reg_data_5; // @[rvdm.scala 393:44:@550.6]
  assign _GEN_56 = _T_168 ? io_dmi_req_bits_data : reg_data_6; // @[rvdm.scala 393:44:@553.6]
  assign _GEN_57 = _T_170 ? io_dmi_req_bits_data : reg_data_7; // @[rvdm.scala 393:44:@556.6]
  assign _GEN_58 = _T_172 ? io_dmi_req_bits_data : reg_data_8; // @[rvdm.scala 393:44:@559.6]
  assign _GEN_59 = _T_174 ? io_dmi_req_bits_data : reg_data_9; // @[rvdm.scala 393:44:@562.6]
  assign _GEN_60 = _T_176 ? io_dmi_req_bits_data : reg_data_10; // @[rvdm.scala 393:44:@565.6]
  assign _GEN_61 = _T_178 ? io_dmi_req_bits_data : reg_data_11; // @[rvdm.scala 393:44:@568.6]
  assign _GEN_63 = _T_384 ? _GEN_21 : reg_abstractcs; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_68 = _T_384 ? _GEN_18 : reg_command; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_69 = _T_384 ? _GEN_19 : reg_regrw; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_75 = _T_384 ? _GEN_27 : reg_dmcontrol; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_81 = _T_384 ? _GEN_33 : reg_sbcs; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_82 = _T_384 ? _GEN_49 : reg_sbaddress_0; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_83 = _T_384 ? _GEN_35 : reg_sbaddress_1; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_84 = _T_384 ? _GEN_36 : reg_sbaddress_2; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_85 = _T_384 ? _GEN_42 : reg_sbdata_0; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_90 = _T_384 ? _GEN_47 : 1'h0; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_91 = _T_384 ? _GEN_48 : 1'h0; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_92 = _T_384 ? _GEN_50 : reg_data_0; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_93 = _T_384 ? _GEN_51 : reg_data_1; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_94 = _T_384 ? _GEN_52 : reg_data_2; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_95 = _T_384 ? _GEN_53 : reg_data_3; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_96 = _T_384 ? _GEN_54 : reg_data_4; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_97 = _T_384 ? _GEN_55 : reg_data_5; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_98 = _T_384 ? _GEN_56 : reg_data_6; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_99 = _T_384 ? _GEN_57 : reg_data_7; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_100 = _T_384 ? _GEN_58 : reg_data_8; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_101 = _T_384 ? _GEN_59 : reg_data_9; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_102 = _T_384 ? _GEN_60 : reg_data_10; // @[rvdm.scala 306:50:@322.4]
  assign _GEN_103 = _T_384 ? _GEN_61 : reg_data_11; // @[rvdm.scala 306:50:@322.4]
  assign _T_514 = 7'h3c == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@578.4]
  assign _T_515 = _T_514 ? reg_sbdata_0 : 32'h0; // @[Mux.scala 46:16:@579.4]
  assign _T_516 = 7'h3b == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@580.4]
  assign _T_517 = _T_516 ? reg_sbaddress_2 : _T_515; // @[Mux.scala 46:16:@581.4]
  assign _T_518 = 7'h3a == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@582.4]
  assign _T_519 = _T_518 ? reg_sbaddress_1 : _T_517; // @[Mux.scala 46:16:@583.4]
  assign _T_520 = 7'h39 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@584.4]
  assign _T_521 = _T_520 ? reg_sbaddress_0 : _T_519; // @[Mux.scala 46:16:@585.4]
  assign _T_522 = 7'h2f == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@586.4]
  assign _T_523 = _T_522 ? 32'h0 : _T_521; // @[Mux.scala 46:16:@587.4]
  assign _T_524 = 7'h2e == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@588.4]
  assign _T_525 = _T_524 ? 32'h0 : _T_523; // @[Mux.scala 46:16:@589.4]
  assign _T_526 = 7'h2d == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@590.4]
  assign _T_527 = _T_526 ? 32'h0 : _T_525; // @[Mux.scala 46:16:@591.4]
  assign _T_528 = 7'h2c == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@592.4]
  assign _T_529 = _T_528 ? 32'h0 : _T_527; // @[Mux.scala 46:16:@593.4]
  assign _T_530 = 7'h2b == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@594.4]
  assign _T_531 = _T_530 ? 32'h0 : _T_529; // @[Mux.scala 46:16:@595.4]
  assign _T_532 = 7'h2a == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@596.4]
  assign _T_533 = _T_532 ? 32'h0 : _T_531; // @[Mux.scala 46:16:@597.4]
  assign _T_534 = 7'h29 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@598.4]
  assign _T_535 = _T_534 ? 32'h0 : _T_533; // @[Mux.scala 46:16:@599.4]
  assign _T_536 = 7'h28 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@600.4]
  assign _T_537 = _T_536 ? 32'h0 : _T_535; // @[Mux.scala 46:16:@601.4]
  assign _T_538 = 7'h27 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@602.4]
  assign _T_539 = _T_538 ? 32'h0 : _T_537; // @[Mux.scala 46:16:@603.4]
  assign _T_540 = 7'h26 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@604.4]
  assign _T_541 = _T_540 ? 32'h0 : _T_539; // @[Mux.scala 46:16:@605.4]
  assign _T_542 = 7'h25 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@606.4]
  assign _T_543 = _T_542 ? 32'h0 : _T_541; // @[Mux.scala 46:16:@607.4]
  assign _T_544 = 7'h24 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@608.4]
  assign _T_545 = _T_544 ? 32'h0 : _T_543; // @[Mux.scala 46:16:@609.4]
  assign _T_546 = 7'h23 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@610.4]
  assign _T_547 = _T_546 ? 32'h0 : _T_545; // @[Mux.scala 46:16:@611.4]
  assign _T_548 = 7'h22 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@612.4]
  assign _T_549 = _T_548 ? 32'h0 : _T_547; // @[Mux.scala 46:16:@613.4]
  assign _T_550 = 7'h21 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@614.4]
  assign _T_551 = _T_550 ? 32'h0 : _T_549; // @[Mux.scala 46:16:@615.4]
  assign _T_552 = 7'h20 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@616.4]
  assign _T_553 = _T_552 ? reg_progbuf_0 : _T_551; // @[Mux.scala 46:16:@617.4]
  assign _T_554 = 7'hf == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@618.4]
  assign _T_555 = _T_554 ? reg_data_11 : _T_553; // @[Mux.scala 46:16:@619.4]
  assign _T_556 = 7'he == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@620.4]
  assign _T_557 = _T_556 ? reg_data_10 : _T_555; // @[Mux.scala 46:16:@621.4]
  assign _T_558 = 7'hd == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@622.4]
  assign _T_559 = _T_558 ? reg_data_9 : _T_557; // @[Mux.scala 46:16:@623.4]
  assign _T_560 = 7'hc == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@624.4]
  assign _T_561 = _T_560 ? reg_data_8 : _T_559; // @[Mux.scala 46:16:@625.4]
  assign _T_562 = 7'hb == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@626.4]
  assign _T_563 = _T_562 ? reg_data_7 : _T_561; // @[Mux.scala 46:16:@627.4]
  assign _T_564 = 7'ha == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@628.4]
  assign _T_565 = _T_564 ? reg_data_6 : _T_563; // @[Mux.scala 46:16:@629.4]
  assign _T_566 = 7'h9 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@630.4]
  assign _T_567 = _T_566 ? reg_data_5 : _T_565; // @[Mux.scala 46:16:@631.4]
  assign _T_568 = 7'h8 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@632.4]
  assign _T_569 = _T_568 ? reg_data_4 : _T_567; // @[Mux.scala 46:16:@633.4]
  assign _T_570 = 7'h7 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@634.4]
  assign _T_571 = _T_570 ? reg_data_3 : _T_569; // @[Mux.scala 46:16:@635.4]
  assign _T_572 = 7'h6 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@636.4]
  assign _T_573 = _T_572 ? reg_data_2 : _T_571; // @[Mux.scala 46:16:@637.4]
  assign _T_574 = 7'h5 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@638.4]
  assign _T_575 = _T_574 ? reg_data_1 : _T_573; // @[Mux.scala 46:16:@639.4]
  assign _T_576 = 7'h4 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@640.4]
  assign _T_577 = _T_576 ? reg_data_0 : _T_575; // @[Mux.scala 46:16:@641.4]
  assign _T_578 = 7'h38 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@642.4]
  assign _T_579 = _T_578 ? reg_sbcs : _T_577; // @[Mux.scala 46:16:@643.4]
  assign _T_580 = 7'h30 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@644.4]
  assign _T_581 = _T_580 ? 32'h0 : _T_579; // @[Mux.scala 46:16:@645.4]
  assign _T_582 = 7'h19 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@646.4]
  assign _T_583 = _T_582 ? 32'h0 : _T_581; // @[Mux.scala 46:16:@647.4]
  assign _T_584 = 7'h18 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@648.4]
  assign _T_585 = _T_584 ? 32'h0 : _T_583; // @[Mux.scala 46:16:@649.4]
  assign _T_586 = 7'h17 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@650.4]
  assign _T_587 = _T_586 ? reg_command : _T_585; // @[Mux.scala 46:16:@651.4]
  assign _T_588 = 7'h16 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@652.4]
  assign _T_589 = _T_588 ? reg_abstractcs : _T_587; // @[Mux.scala 46:16:@653.4]
  assign _T_590 = 7'h15 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@654.4]
  assign _T_591 = _T_590 ? 32'h0 : _T_589; // @[Mux.scala 46:16:@655.4]
  assign _T_592 = 7'h14 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@656.4]
  assign _T_593 = _T_592 ? 32'h0 : _T_591; // @[Mux.scala 46:16:@657.4]
  assign _T_594 = 7'h13 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@658.4]
  assign _T_595 = _T_594 ? 32'h0 : _T_593; // @[Mux.scala 46:16:@659.4]
  assign _T_596 = 7'h12 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@660.4]
  assign _T_597 = _T_596 ? 32'h111bc0 : _T_595; // @[Mux.scala 46:16:@661.4]
  assign _T_598 = 7'h11 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@662.4]
  assign _T_599 = _T_598 ? reg_dmstatus : _T_597; // @[Mux.scala 46:16:@663.4]
  assign _T_600 = 7'h10 == io_dmi_req_bits_addr; // @[Mux.scala 46:19:@664.4]
  assign _T_601 = _T_600 ? reg_dmcontrol : _T_599; // @[Mux.scala 46:16:@665.4]
  assign _T_604 = command_regno & 16'h1f; // @[rvdm.scala 404:38:@668.4]
  assign _T_605 = _T_604[4:0]; // @[rvdm.scala 404:47:@669.4]
  assign cmd_regrw = command_transfer & reg_regrw; // @[rvdm.scala 406:39:@671.4]
  assign _GEN_106 = command_write ? _GEN_92 : io_ddpath_rdata; // @[rvdm.scala 408:29:@673.6]
  assign _GEN_108 = cmd_regrw ? command_write : 1'h0; // @[rvdm.scala 407:21:@672.4]
  assign _GEN_109 = cmd_regrw ? _GEN_106 : _GEN_92; // @[rvdm.scala 407:21:@672.4]
  assign _GEN_110 = cmd_regrw ? 1'h0 : _GEN_69; // @[rvdm.scala 407:21:@672.4]
  assign _T_608 = io_dmi_req_bits_op == 2'h1; // @[rvdm.scala 424:29:@682.4]
  assign _T_609 = _T_608 & _T_218; // @[rvdm.scala 424:47:@683.4]
  assign _T_611 = io_ddmem_resp_valid & reg_ddmem_req_valid; // @[rvdm.scala 434:37:@690.8]
  assign _GEN_111 = sbcs_sbautoincrement ? _T_506 : _GEN_82; // @[rvdm.scala 441:44:@696.10]
  assign _GEN_113 = _T_611 ? io_ddmem_resp_data : _GEN_85; // @[rvdm.scala 434:59:@691.8]
  assign _GEN_114 = _T_611 ? 1'h0 : 1'h1; // @[rvdm.scala 434:59:@691.8]
  assign _GEN_115 = _T_611 ? 1'h0 : reg_mrdata_requested; // @[rvdm.scala 434:59:@691.8]
  assign _GEN_116 = _T_611 ? 1'h1 : _GEN_91; // @[rvdm.scala 434:59:@691.8]
  assign _GEN_117 = _T_611 ? _GEN_111 : _GEN_82; // @[rvdm.scala 434:59:@691.8]
  assign _GEN_118 = io_ddmem_req_ready ? 1'h1 : reg_mrdata_requested; // @[rvdm.scala 455:38:@711.8]
  assign _GEN_119 = reg_mrdata_requested ? _GEN_114 : _GEN_37; // @[rvdm.scala 432:36:@688.6]
  assign _GEN_120 = reg_mrdata_requested ? _GEN_113 : _GEN_85; // @[rvdm.scala 432:36:@688.6]
  assign _GEN_121 = reg_mrdata_requested ? _GEN_115 : _GEN_118; // @[rvdm.scala 432:36:@688.6]
  assign _GEN_122 = reg_mrdata_requested ? _GEN_116 : _GEN_91; // @[rvdm.scala 432:36:@688.6]
  assign _GEN_123 = reg_mrdata_requested ? _GEN_117 : _GEN_82; // @[rvdm.scala 432:36:@688.6]
  assign _GEN_124 = _T_609 ? 1'h0 : 1'h1; // @[rvdm.scala 424:74:@684.4]
  assign _GEN_127 = _T_609 ? _GEN_119 : _GEN_90; // @[rvdm.scala 424:74:@684.4]
  assign _GEN_128 = _T_609 ? _GEN_120 : _GEN_85; // @[rvdm.scala 424:74:@684.4]
  assign _GEN_129 = _T_609 ? _GEN_121 : reg_mrdata_requested; // @[rvdm.scala 424:74:@684.4]
  assign _GEN_130 = _T_609 ? _GEN_122 : _GEN_91; // @[rvdm.scala 424:74:@684.4]
  assign _GEN_131 = _T_609 ? _GEN_123 : _GEN_82; // @[rvdm.scala 424:74:@684.4]
  assign _T_623 = _T_218 == 1'h0; // @[rvdm.scala 463:10:@716.4]
  assign _GEN_132 = _T_623 ? 1'h0 : _GEN_129; // @[rvdm.scala 463:39:@717.4]
  assign _T_625 = _T_218 ? reg_delay_mrwdata_valid : io_dmi_req_ready; // @[rvdm.scala 479:29:@720.4]
  assign _T_627 = io_dmi_req_bits_addr == 7'h44; // @[rvdm.scala 490:32:@724.4]
  assign _T_628 = _T_627 & io_dmi_req_valid; // @[rvdm.scala 490:45:@725.4]
  assign _GEN_133 = _T_628 ? 1'h0 : reg_rstcore; // @[rvdm.scala 490:65:@726.4]
  assign _T_631 = io_dmi_req_bits_addr == 7'h48; // @[rvdm.scala 493:32:@729.4]
  assign _T_632 = _T_631 & io_dmi_req_valid; // @[rvdm.scala 493:45:@730.4]
  assign _GEN_134 = _T_632 ? 1'h1 : _GEN_133; // @[rvdm.scala 493:65:@731.4]
  assign _GEN_135 = reset ? 32'h0 : _GEN_75; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_136 = reset ? _T_498 : _GEN_81; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_137 = reset ? 32'h0 : _GEN_68; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_138 = reset ? 32'h0 : reg_progbuf_0; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_139 = reset ? 32'h0 : _GEN_109; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_140 = reset ? 32'h0 : _GEN_131; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_141 = reset ? 32'h0 : _GEN_128; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_142 = reset ? 1'h0 : _GEN_127; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_143 = reset ? 1'h0 : _GEN_108; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_146 = reset ? _T_380 : _T_380; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_152 = reset ? _T_404 : _GEN_63; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_153 = reset ? 1'h0 : _GEN_132; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_154 = reset ? 1'h0 : _GEN_130; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_155 = reset ? 2'h3 : 2'h0; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_156 = reset ? 1'h0 : _GEN_110; // @[rvdm.scala 498:26:@735.4]
  assign _GEN_157 = reset ? 1'h1 : _GEN_134; // @[rvdm.scala 498:26:@735.4]
  assign io_dmi_req_ready = io_dmi_req_valid;
  assign io_dmi_resp_bits_resp = _GEN_155;
  assign io_dmi_resp_bits_data = _T_601;
  assign io_dmi_resp_valid = _T_625;
  assign io_ddpath_addr = _T_605;
  assign io_ddpath_wdata = reg_data_0;
  assign io_ddpath_valid = _GEN_143;
  assign io_ddmem_req_addr = reg_sbaddress_0;
  assign io_ddmem_req_data = reg_sbdata_0;
  assign io_ddmem_req_mfunc = _GEN_124;
  assign io_ddmem_req_valid = reg_ddmem_req_valid;
  assign io_rstcore = reg_rstcore;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  reg_dmstatus = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  reg_dmcontrol = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  reg_sbcs = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  reg_abstractcs = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  reg_command = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  reg_progbuf_0 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  reg_data_0 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  reg_data_1 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  reg_data_2 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  reg_data_3 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  reg_data_4 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  reg_data_5 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  reg_data_6 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  reg_data_7 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  reg_data_8 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  reg_data_9 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  reg_data_10 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  reg_data_11 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  reg_sbaddress_0 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  reg_sbaddress_1 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  reg_sbaddress_2 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  reg_sbdata_0 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  reg_regrw = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  reg_mrdata_requested = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  reg_delay_mrwdata_valid = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  reg_ddmem_req_valid = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  reg_rstcore = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    reg_dmstatus <= {{2'd0}, _GEN_146};
    if (reset) begin
      reg_dmcontrol <= 32'h0;
    end else begin
      if (_T_384) begin
        if (_T_132) begin
          reg_dmcontrol <= _T_470;
        end
      end
    end
    if (reset) begin
      reg_sbcs <= _T_498;
    end else begin
      if (_T_384) begin
        if (_T_154) begin
          reg_sbcs <= _T_498;
        end
      end
    end
    if (reset) begin
      reg_abstractcs <= _T_404;
    end else begin
      if (_T_384) begin
        if (_T_146) begin
          if (_T_419) begin
            reg_abstractcs <= _T_404;
          end else begin
            reg_abstractcs <= _T_404;
          end
        end else begin
          if (_T_144) begin
            if (io_dmi_req_valid) begin
              reg_abstractcs <= _T_404;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_command <= 32'h0;
    end else begin
      if (_T_384) begin
        if (_T_146) begin
          if (_T_419) begin
            reg_command <= _T_426;
          end
        end
      end
    end
    if (reset) begin
      reg_progbuf_0 <= 32'h0;
    end
    if (reset) begin
      reg_data_0 <= 32'h0;
    end else begin
      if (cmd_regrw) begin
        if (command_write) begin
          if (_T_384) begin
            if (_T_156) begin
              reg_data_0 <= io_dmi_req_bits_data;
            end
          end
        end else begin
          reg_data_0 <= io_ddpath_rdata;
        end
      end else begin
        if (_T_384) begin
          if (_T_156) begin
            reg_data_0 <= io_dmi_req_bits_data;
          end
        end
      end
    end
    if (_T_384) begin
      if (_T_158) begin
        reg_data_1 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_160) begin
        reg_data_2 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_162) begin
        reg_data_3 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_164) begin
        reg_data_4 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_166) begin
        reg_data_5 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_168) begin
        reg_data_6 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_170) begin
        reg_data_7 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_172) begin
        reg_data_8 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_174) begin
        reg_data_9 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_176) begin
        reg_data_10 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_178) begin
        reg_data_11 <= io_dmi_req_bits_data;
      end
    end
    if (reset) begin
      reg_sbaddress_0 <= 32'h0;
    end else begin
      if (_T_609) begin
        if (reg_mrdata_requested) begin
          if (_T_611) begin
            if (sbcs_sbautoincrement) begin
              reg_sbaddress_0 <= _T_506;
            end else begin
              if (_T_384) begin
                if (_T_218) begin
                  if (_T_501) begin
                    if (sbcs_sbautoincrement) begin
                      reg_sbaddress_0 <= _T_506;
                    end else begin
                      if (_T_212) begin
                        reg_sbaddress_0 <= io_dmi_req_bits_data;
                      end
                    end
                  end else begin
                    if (_T_212) begin
                      reg_sbaddress_0 <= io_dmi_req_bits_data;
                    end
                  end
                end else begin
                  if (_T_212) begin
                    reg_sbaddress_0 <= io_dmi_req_bits_data;
                  end
                end
              end
            end
          end else begin
            if (_T_384) begin
              if (_T_218) begin
                if (_T_501) begin
                  if (sbcs_sbautoincrement) begin
                    reg_sbaddress_0 <= _T_506;
                  end else begin
                    if (_T_212) begin
                      reg_sbaddress_0 <= io_dmi_req_bits_data;
                    end
                  end
                end else begin
                  reg_sbaddress_0 <= _GEN_34;
                end
              end else begin
                reg_sbaddress_0 <= _GEN_34;
              end
            end
          end
        end else begin
          if (_T_384) begin
            if (_T_218) begin
              if (_T_501) begin
                if (sbcs_sbautoincrement) begin
                  reg_sbaddress_0 <= _T_506;
                end else begin
                  reg_sbaddress_0 <= _GEN_34;
                end
              end else begin
                reg_sbaddress_0 <= _GEN_34;
              end
            end else begin
              reg_sbaddress_0 <= _GEN_34;
            end
          end
        end
      end else begin
        if (_T_384) begin
          if (_T_218) begin
            if (_T_501) begin
              if (sbcs_sbautoincrement) begin
                reg_sbaddress_0 <= _T_506;
              end else begin
                reg_sbaddress_0 <= _GEN_34;
              end
            end else begin
              reg_sbaddress_0 <= _GEN_34;
            end
          end else begin
            reg_sbaddress_0 <= _GEN_34;
          end
        end
      end
    end
    if (_T_384) begin
      if (_T_214) begin
        reg_sbaddress_1 <= io_dmi_req_bits_data;
      end
    end
    if (_T_384) begin
      if (_T_216) begin
        reg_sbaddress_2 <= io_dmi_req_bits_data;
      end
    end
    if (reset) begin
      reg_sbdata_0 <= 32'h0;
    end else begin
      if (_T_609) begin
        if (reg_mrdata_requested) begin
          if (_T_611) begin
            reg_sbdata_0 <= io_ddmem_resp_data;
          end else begin
            if (_T_384) begin
              if (_T_218) begin
                reg_sbdata_0 <= io_dmi_req_bits_data;
              end
            end
          end
        end else begin
          if (_T_384) begin
            if (_T_218) begin
              reg_sbdata_0 <= io_dmi_req_bits_data;
            end
          end
        end
      end else begin
        if (_T_384) begin
          if (_T_218) begin
            reg_sbdata_0 <= io_dmi_req_bits_data;
          end
        end
      end
    end
    if (reset) begin
      reg_regrw <= 1'h0;
    end else begin
      if (cmd_regrw) begin
        reg_regrw <= 1'h0;
      end else begin
        if (_T_384) begin
          if (_T_146) begin
            if (_T_419) begin
              reg_regrw <= _T_412;
            end else begin
              reg_regrw <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mrdata_requested <= 1'h0;
    end else begin
      if (_T_623) begin
        reg_mrdata_requested <= 1'h0;
      end else begin
        if (_T_609) begin
          if (reg_mrdata_requested) begin
            if (_T_611) begin
              reg_mrdata_requested <= 1'h0;
            end
          end else begin
            if (io_ddmem_req_ready) begin
              reg_mrdata_requested <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_delay_mrwdata_valid <= 1'h0;
    end else begin
      if (_T_609) begin
        if (reg_mrdata_requested) begin
          if (_T_611) begin
            reg_delay_mrwdata_valid <= 1'h1;
          end else begin
            if (_T_384) begin
              if (_T_218) begin
                reg_delay_mrwdata_valid <= _T_501;
              end else begin
                reg_delay_mrwdata_valid <= 1'h0;
              end
            end else begin
              reg_delay_mrwdata_valid <= 1'h0;
            end
          end
        end else begin
          if (_T_384) begin
            if (_T_218) begin
              reg_delay_mrwdata_valid <= _T_501;
            end else begin
              reg_delay_mrwdata_valid <= 1'h0;
            end
          end else begin
            reg_delay_mrwdata_valid <= 1'h0;
          end
        end
      end else begin
        if (_T_384) begin
          if (_T_218) begin
            reg_delay_mrwdata_valid <= _T_501;
          end else begin
            reg_delay_mrwdata_valid <= 1'h0;
          end
        end else begin
          reg_delay_mrwdata_valid <= 1'h0;
        end
      end
    end
    if (reset) begin
      reg_ddmem_req_valid <= 1'h0;
    end else begin
      if (_T_609) begin
        if (reg_mrdata_requested) begin
          if (_T_611) begin
            reg_ddmem_req_valid <= 1'h0;
          end else begin
            reg_ddmem_req_valid <= 1'h1;
          end
        end else begin
          if (reg_delay_mrwdata_valid) begin
            reg_ddmem_req_valid <= 1'h0;
          end else begin
            reg_ddmem_req_valid <= 1'h1;
          end
        end
      end else begin
        if (_T_384) begin
          if (_T_218) begin
            if (_T_501) begin
              reg_ddmem_req_valid <= 1'h0;
            end else begin
              if (reg_delay_mrwdata_valid) begin
                reg_ddmem_req_valid <= 1'h0;
              end else begin
                reg_ddmem_req_valid <= 1'h1;
              end
            end
          end else begin
            reg_ddmem_req_valid <= 1'h0;
          end
        end else begin
          reg_ddmem_req_valid <= 1'h0;
        end
      end
    end
    if (reset) begin
      reg_rstcore <= 1'h1;
    end else begin
      if (_T_632) begin
        reg_rstcore <= 1'h1;
      end else begin
        if (_T_628) begin
          reg_rstcore <= 1'h0;
        end
      end
    end
  end
endmodule
module rvcpath( // @[:@800.2]
  input  [31:0] io_d2c_inst, // @[:@803.4]
  input         io_d2c_dexcp, // @[:@803.4]
  output [3:0]  io_c2d_alu_func, // @[:@803.4]
  output [2:0]  io_c2d_op2_sel, // @[:@803.4]
  output        io_c2d_reg_wren, // @[:@803.4]
  output        io_c2d_mem_wren, // @[:@803.4]
  output        io_c2d_mem_en, // @[:@803.4]
  output [1:0]  io_c2d_wb_sel, // @[:@803.4]
  output [2:0]  io_c2d_mem_type, // @[:@803.4]
  output [1:0]  io_c2d_pc_sel, // @[:@803.4]
  output [2:0]  io_c2d_br_sel, // @[:@803.4]
  output [1:0]  io_c2d_op1_sel, // @[:@803.4]
  output [2:0]  io_c2d_csr_cmd, // @[:@803.4]
  output        io_c2d_cexcp, // @[:@803.4]
  output [3:0]  io_c2d_ccause // @[:@803.4]
);
  wire [31:0] _T_123; // @[Lookup.scala 9:38:@837.4]
  wire  _T_124; // @[Lookup.scala 9:38:@838.4]
  wire  _T_128; // @[Lookup.scala 9:38:@840.4]
  wire  _T_132; // @[Lookup.scala 9:38:@842.4]
  wire [31:0] _T_135; // @[Lookup.scala 9:38:@843.4]
  wire  _T_136; // @[Lookup.scala 9:38:@844.4]
  wire  _T_140; // @[Lookup.scala 9:38:@846.4]
  wire  _T_144; // @[Lookup.scala 9:38:@848.4]
  wire  _T_148; // @[Lookup.scala 9:38:@850.4]
  wire  _T_152; // @[Lookup.scala 9:38:@852.4]
  wire  _T_156; // @[Lookup.scala 9:38:@854.4]
  wire  _T_160; // @[Lookup.scala 9:38:@856.4]
  wire  _T_164; // @[Lookup.scala 9:38:@858.4]
  wire  _T_168; // @[Lookup.scala 9:38:@860.4]
  wire  _T_172; // @[Lookup.scala 9:38:@862.4]
  wire  _T_176; // @[Lookup.scala 9:38:@864.4]
  wire  _T_180; // @[Lookup.scala 9:38:@866.4]
  wire  _T_184; // @[Lookup.scala 9:38:@868.4]
  wire  _T_188; // @[Lookup.scala 9:38:@870.4]
  wire  _T_192; // @[Lookup.scala 9:38:@872.4]
  wire  _T_196; // @[Lookup.scala 9:38:@874.4]
  wire  _T_200; // @[Lookup.scala 9:38:@876.4]
  wire  _T_204; // @[Lookup.scala 9:38:@878.4]
  wire  _T_208; // @[Lookup.scala 9:38:@880.4]
  wire  _T_212; // @[Lookup.scala 9:38:@882.4]
  wire  _T_216; // @[Lookup.scala 9:38:@884.4]
  wire [31:0] _T_219; // @[Lookup.scala 9:38:@885.4]
  wire  _T_220; // @[Lookup.scala 9:38:@886.4]
  wire  _T_224; // @[Lookup.scala 9:38:@888.4]
  wire  _T_228; // @[Lookup.scala 9:38:@890.4]
  wire  _T_232; // @[Lookup.scala 9:38:@892.4]
  wire  _T_236; // @[Lookup.scala 9:38:@894.4]
  wire  _T_240; // @[Lookup.scala 9:38:@896.4]
  wire  _T_244; // @[Lookup.scala 9:38:@898.4]
  wire  _T_248; // @[Lookup.scala 9:38:@900.4]
  wire  _T_252; // @[Lookup.scala 9:38:@902.4]
  wire  _T_256; // @[Lookup.scala 9:38:@904.4]
  wire  _T_260; // @[Lookup.scala 9:38:@906.4]
  wire  _T_264; // @[Lookup.scala 9:38:@908.4]
  wire  _T_268; // @[Lookup.scala 9:38:@910.4]
  wire  _T_272; // @[Lookup.scala 9:38:@912.4]
  wire  _T_276; // @[Lookup.scala 9:38:@914.4]
  wire  _T_280; // @[Lookup.scala 9:38:@916.4]
  wire  _T_284; // @[Lookup.scala 9:38:@918.4]
  wire  _T_288; // @[Lookup.scala 9:38:@920.4]
  wire  _T_292; // @[Lookup.scala 9:38:@922.4]
  wire [31:0] _T_295; // @[Lookup.scala 9:38:@923.4]
  wire  _T_296; // @[Lookup.scala 9:38:@924.4]
  wire  _T_300; // @[Lookup.scala 9:38:@926.4]
  wire  _T_304; // @[Lookup.scala 9:38:@928.4]
  wire  _T_308; // @[Lookup.scala 9:38:@930.4]
  wire  _T_312; // @[Lookup.scala 9:38:@932.4]
  wire  _T_316; // @[Lookup.scala 9:38:@934.4]
  wire  _T_320; // @[Lookup.scala 9:38:@936.4]
  wire [3:0] _T_334; // @[Lookup.scala 11:37:@950.4]
  wire [3:0] _T_335; // @[Lookup.scala 11:37:@951.4]
  wire [3:0] _T_336; // @[Lookup.scala 11:37:@952.4]
  wire [3:0] _T_337; // @[Lookup.scala 11:37:@953.4]
  wire [3:0] _T_338; // @[Lookup.scala 11:37:@954.4]
  wire [3:0] _T_339; // @[Lookup.scala 11:37:@955.4]
  wire [3:0] _T_340; // @[Lookup.scala 11:37:@956.4]
  wire [3:0] _T_341; // @[Lookup.scala 11:37:@957.4]
  wire [3:0] _T_342; // @[Lookup.scala 11:37:@958.4]
  wire [3:0] _T_343; // @[Lookup.scala 11:37:@959.4]
  wire [3:0] _T_344; // @[Lookup.scala 11:37:@960.4]
  wire [3:0] _T_345; // @[Lookup.scala 11:37:@961.4]
  wire [3:0] _T_346; // @[Lookup.scala 11:37:@962.4]
  wire [3:0] _T_347; // @[Lookup.scala 11:37:@963.4]
  wire [3:0] _T_348; // @[Lookup.scala 11:37:@964.4]
  wire [3:0] _T_349; // @[Lookup.scala 11:37:@965.4]
  wire [3:0] _T_350; // @[Lookup.scala 11:37:@966.4]
  wire [3:0] _T_351; // @[Lookup.scala 11:37:@967.4]
  wire [3:0] _T_352; // @[Lookup.scala 11:37:@968.4]
  wire [3:0] _T_353; // @[Lookup.scala 11:37:@969.4]
  wire [3:0] _T_354; // @[Lookup.scala 11:37:@970.4]
  wire [3:0] _T_355; // @[Lookup.scala 11:37:@971.4]
  wire [3:0] _T_356; // @[Lookup.scala 11:37:@972.4]
  wire [3:0] _T_357; // @[Lookup.scala 11:37:@973.4]
  wire [3:0] _T_358; // @[Lookup.scala 11:37:@974.4]
  wire [3:0] _T_359; // @[Lookup.scala 11:37:@975.4]
  wire [3:0] _T_360; // @[Lookup.scala 11:37:@976.4]
  wire [3:0] _T_361; // @[Lookup.scala 11:37:@977.4]
  wire [3:0] _T_362; // @[Lookup.scala 11:37:@978.4]
  wire [3:0] _T_363; // @[Lookup.scala 11:37:@979.4]
  wire [3:0] _T_364; // @[Lookup.scala 11:37:@980.4]
  wire [3:0] _T_365; // @[Lookup.scala 11:37:@981.4]
  wire [3:0] _T_366; // @[Lookup.scala 11:37:@982.4]
  wire [3:0] _T_367; // @[Lookup.scala 11:37:@983.4]
  wire [3:0] _T_368; // @[Lookup.scala 11:37:@984.4]
  wire [3:0] _T_369; // @[Lookup.scala 11:37:@985.4]
  wire [3:0] alu_func; // @[Lookup.scala 11:37:@986.4]
  wire [2:0] _T_383; // @[Lookup.scala 11:37:@1000.4]
  wire [2:0] _T_384; // @[Lookup.scala 11:37:@1001.4]
  wire [2:0] _T_385; // @[Lookup.scala 11:37:@1002.4]
  wire [2:0] _T_386; // @[Lookup.scala 11:37:@1003.4]
  wire [2:0] _T_387; // @[Lookup.scala 11:37:@1004.4]
  wire [2:0] _T_388; // @[Lookup.scala 11:37:@1005.4]
  wire [2:0] _T_389; // @[Lookup.scala 11:37:@1006.4]
  wire [2:0] _T_390; // @[Lookup.scala 11:37:@1007.4]
  wire [2:0] _T_391; // @[Lookup.scala 11:37:@1008.4]
  wire [2:0] _T_392; // @[Lookup.scala 11:37:@1009.4]
  wire [2:0] _T_393; // @[Lookup.scala 11:37:@1010.4]
  wire [2:0] _T_394; // @[Lookup.scala 11:37:@1011.4]
  wire [2:0] _T_395; // @[Lookup.scala 11:37:@1012.4]
  wire [2:0] _T_396; // @[Lookup.scala 11:37:@1013.4]
  wire [2:0] _T_397; // @[Lookup.scala 11:37:@1014.4]
  wire [2:0] _T_398; // @[Lookup.scala 11:37:@1015.4]
  wire [2:0] _T_399; // @[Lookup.scala 11:37:@1016.4]
  wire [2:0] _T_400; // @[Lookup.scala 11:37:@1017.4]
  wire [2:0] _T_401; // @[Lookup.scala 11:37:@1018.4]
  wire [2:0] _T_402; // @[Lookup.scala 11:37:@1019.4]
  wire [2:0] _T_403; // @[Lookup.scala 11:37:@1020.4]
  wire [2:0] _T_404; // @[Lookup.scala 11:37:@1021.4]
  wire [2:0] _T_405; // @[Lookup.scala 11:37:@1022.4]
  wire [2:0] _T_406; // @[Lookup.scala 11:37:@1023.4]
  wire [2:0] _T_407; // @[Lookup.scala 11:37:@1024.4]
  wire [2:0] _T_408; // @[Lookup.scala 11:37:@1025.4]
  wire [2:0] _T_409; // @[Lookup.scala 11:37:@1026.4]
  wire [2:0] _T_410; // @[Lookup.scala 11:37:@1027.4]
  wire [2:0] _T_411; // @[Lookup.scala 11:37:@1028.4]
  wire [2:0] _T_412; // @[Lookup.scala 11:37:@1029.4]
  wire [2:0] _T_413; // @[Lookup.scala 11:37:@1030.4]
  wire [2:0] _T_414; // @[Lookup.scala 11:37:@1031.4]
  wire [2:0] _T_415; // @[Lookup.scala 11:37:@1032.4]
  wire [2:0] _T_416; // @[Lookup.scala 11:37:@1033.4]
  wire [2:0] _T_417; // @[Lookup.scala 11:37:@1034.4]
  wire [2:0] _T_418; // @[Lookup.scala 11:37:@1035.4]
  wire [2:0] ctlsig_1; // @[Lookup.scala 11:37:@1036.4]
  wire  _T_427; // @[Lookup.scala 11:37:@1045.4]
  wire  _T_428; // @[Lookup.scala 11:37:@1046.4]
  wire  _T_429; // @[Lookup.scala 11:37:@1047.4]
  wire  _T_430; // @[Lookup.scala 11:37:@1048.4]
  wire  _T_431; // @[Lookup.scala 11:37:@1049.4]
  wire  _T_432; // @[Lookup.scala 11:37:@1050.4]
  wire  _T_433; // @[Lookup.scala 11:37:@1051.4]
  wire  _T_434; // @[Lookup.scala 11:37:@1052.4]
  wire  _T_435; // @[Lookup.scala 11:37:@1053.4]
  wire  _T_436; // @[Lookup.scala 11:37:@1054.4]
  wire  _T_437; // @[Lookup.scala 11:37:@1055.4]
  wire  _T_438; // @[Lookup.scala 11:37:@1056.4]
  wire  _T_439; // @[Lookup.scala 11:37:@1057.4]
  wire  _T_440; // @[Lookup.scala 11:37:@1058.4]
  wire  _T_441; // @[Lookup.scala 11:37:@1059.4]
  wire  _T_442; // @[Lookup.scala 11:37:@1060.4]
  wire  _T_443; // @[Lookup.scala 11:37:@1061.4]
  wire  _T_444; // @[Lookup.scala 11:37:@1062.4]
  wire  _T_445; // @[Lookup.scala 11:37:@1063.4]
  wire  _T_446; // @[Lookup.scala 11:37:@1064.4]
  wire  _T_447; // @[Lookup.scala 11:37:@1065.4]
  wire  _T_448; // @[Lookup.scala 11:37:@1066.4]
  wire  _T_449; // @[Lookup.scala 11:37:@1067.4]
  wire  _T_450; // @[Lookup.scala 11:37:@1068.4]
  wire  _T_451; // @[Lookup.scala 11:37:@1069.4]
  wire  _T_452; // @[Lookup.scala 11:37:@1070.4]
  wire  _T_453; // @[Lookup.scala 11:37:@1071.4]
  wire  _T_454; // @[Lookup.scala 11:37:@1072.4]
  wire  _T_455; // @[Lookup.scala 11:37:@1073.4]
  wire  _T_456; // @[Lookup.scala 11:37:@1074.4]
  wire  _T_457; // @[Lookup.scala 11:37:@1075.4]
  wire  _T_458; // @[Lookup.scala 11:37:@1076.4]
  wire  _T_459; // @[Lookup.scala 11:37:@1077.4]
  wire  _T_460; // @[Lookup.scala 11:37:@1078.4]
  wire  _T_461; // @[Lookup.scala 11:37:@1079.4]
  wire  _T_462; // @[Lookup.scala 11:37:@1080.4]
  wire  _T_463; // @[Lookup.scala 11:37:@1081.4]
  wire  _T_464; // @[Lookup.scala 11:37:@1082.4]
  wire  _T_465; // @[Lookup.scala 11:37:@1083.4]
  wire  _T_466; // @[Lookup.scala 11:37:@1084.4]
  wire  _T_467; // @[Lookup.scala 11:37:@1085.4]
  wire  ctlsig_2; // @[Lookup.scala 11:37:@1086.4]
  wire  _T_501; // @[Lookup.scala 11:37:@1120.4]
  wire  _T_502; // @[Lookup.scala 11:37:@1121.4]
  wire  _T_503; // @[Lookup.scala 11:37:@1122.4]
  wire  _T_504; // @[Lookup.scala 11:37:@1123.4]
  wire  _T_505; // @[Lookup.scala 11:37:@1124.4]
  wire  _T_506; // @[Lookup.scala 11:37:@1125.4]
  wire  _T_507; // @[Lookup.scala 11:37:@1126.4]
  wire  _T_508; // @[Lookup.scala 11:37:@1127.4]
  wire  _T_509; // @[Lookup.scala 11:37:@1128.4]
  wire  _T_510; // @[Lookup.scala 11:37:@1129.4]
  wire  _T_511; // @[Lookup.scala 11:37:@1130.4]
  wire  _T_512; // @[Lookup.scala 11:37:@1131.4]
  wire  _T_513; // @[Lookup.scala 11:37:@1132.4]
  wire  _T_514; // @[Lookup.scala 11:37:@1133.4]
  wire  _T_515; // @[Lookup.scala 11:37:@1134.4]
  wire  _T_516; // @[Lookup.scala 11:37:@1135.4]
  wire  ctlsig_3; // @[Lookup.scala 11:37:@1136.4]
  wire  _T_552; // @[Lookup.scala 11:37:@1172.4]
  wire  _T_553; // @[Lookup.scala 11:37:@1173.4]
  wire  _T_554; // @[Lookup.scala 11:37:@1174.4]
  wire  _T_555; // @[Lookup.scala 11:37:@1175.4]
  wire  _T_556; // @[Lookup.scala 11:37:@1176.4]
  wire  _T_557; // @[Lookup.scala 11:37:@1177.4]
  wire  _T_558; // @[Lookup.scala 11:37:@1178.4]
  wire  _T_559; // @[Lookup.scala 11:37:@1179.4]
  wire  _T_560; // @[Lookup.scala 11:37:@1180.4]
  wire  _T_561; // @[Lookup.scala 11:37:@1181.4]
  wire  _T_562; // @[Lookup.scala 11:37:@1182.4]
  wire  _T_563; // @[Lookup.scala 11:37:@1183.4]
  wire  _T_564; // @[Lookup.scala 11:37:@1184.4]
  wire  _T_565; // @[Lookup.scala 11:37:@1185.4]
  wire  ctlsig_4; // @[Lookup.scala 11:37:@1186.4]
  wire [1:0] _T_573; // @[Lookup.scala 11:37:@1194.4]
  wire [1:0] _T_574; // @[Lookup.scala 11:37:@1195.4]
  wire [1:0] _T_575; // @[Lookup.scala 11:37:@1196.4]
  wire [1:0] _T_576; // @[Lookup.scala 11:37:@1197.4]
  wire [1:0] _T_577; // @[Lookup.scala 11:37:@1198.4]
  wire [1:0] _T_578; // @[Lookup.scala 11:37:@1199.4]
  wire [1:0] _T_579; // @[Lookup.scala 11:37:@1200.4]
  wire [1:0] _T_580; // @[Lookup.scala 11:37:@1201.4]
  wire [1:0] _T_581; // @[Lookup.scala 11:37:@1202.4]
  wire [1:0] _T_582; // @[Lookup.scala 11:37:@1203.4]
  wire [1:0] _T_583; // @[Lookup.scala 11:37:@1204.4]
  wire [1:0] _T_584; // @[Lookup.scala 11:37:@1205.4]
  wire [1:0] _T_585; // @[Lookup.scala 11:37:@1206.4]
  wire [1:0] _T_586; // @[Lookup.scala 11:37:@1207.4]
  wire [1:0] _T_587; // @[Lookup.scala 11:37:@1208.4]
  wire [1:0] _T_588; // @[Lookup.scala 11:37:@1209.4]
  wire [1:0] _T_589; // @[Lookup.scala 11:37:@1210.4]
  wire [1:0] _T_590; // @[Lookup.scala 11:37:@1211.4]
  wire [1:0] _T_591; // @[Lookup.scala 11:37:@1212.4]
  wire [1:0] _T_592; // @[Lookup.scala 11:37:@1213.4]
  wire [1:0] _T_593; // @[Lookup.scala 11:37:@1214.4]
  wire [1:0] _T_594; // @[Lookup.scala 11:37:@1215.4]
  wire [1:0] _T_595; // @[Lookup.scala 11:37:@1216.4]
  wire [1:0] _T_596; // @[Lookup.scala 11:37:@1217.4]
  wire [1:0] _T_597; // @[Lookup.scala 11:37:@1218.4]
  wire [1:0] _T_598; // @[Lookup.scala 11:37:@1219.4]
  wire [1:0] _T_599; // @[Lookup.scala 11:37:@1220.4]
  wire [1:0] _T_600; // @[Lookup.scala 11:37:@1221.4]
  wire [1:0] _T_601; // @[Lookup.scala 11:37:@1222.4]
  wire [1:0] _T_602; // @[Lookup.scala 11:37:@1223.4]
  wire [1:0] _T_603; // @[Lookup.scala 11:37:@1224.4]
  wire [1:0] _T_604; // @[Lookup.scala 11:37:@1225.4]
  wire [1:0] _T_605; // @[Lookup.scala 11:37:@1226.4]
  wire [1:0] _T_606; // @[Lookup.scala 11:37:@1227.4]
  wire [1:0] _T_607; // @[Lookup.scala 11:37:@1228.4]
  wire [1:0] _T_608; // @[Lookup.scala 11:37:@1229.4]
  wire [1:0] _T_609; // @[Lookup.scala 11:37:@1230.4]
  wire [1:0] _T_610; // @[Lookup.scala 11:37:@1231.4]
  wire [1:0] _T_611; // @[Lookup.scala 11:37:@1232.4]
  wire [1:0] _T_612; // @[Lookup.scala 11:37:@1233.4]
  wire [1:0] _T_613; // @[Lookup.scala 11:37:@1234.4]
  wire [1:0] _T_614; // @[Lookup.scala 11:37:@1235.4]
  wire [1:0] ctlsig_5; // @[Lookup.scala 11:37:@1236.4]
  wire [2:0] _T_648; // @[Lookup.scala 11:37:@1270.4]
  wire [2:0] _T_649; // @[Lookup.scala 11:37:@1271.4]
  wire [2:0] _T_650; // @[Lookup.scala 11:37:@1272.4]
  wire [2:0] _T_651; // @[Lookup.scala 11:37:@1273.4]
  wire [2:0] _T_652; // @[Lookup.scala 11:37:@1274.4]
  wire [2:0] _T_653; // @[Lookup.scala 11:37:@1275.4]
  wire [2:0] _T_654; // @[Lookup.scala 11:37:@1276.4]
  wire [2:0] _T_655; // @[Lookup.scala 11:37:@1277.4]
  wire [2:0] _T_656; // @[Lookup.scala 11:37:@1278.4]
  wire [2:0] _T_657; // @[Lookup.scala 11:37:@1279.4]
  wire [2:0] _T_658; // @[Lookup.scala 11:37:@1280.4]
  wire [2:0] _T_659; // @[Lookup.scala 11:37:@1281.4]
  wire [2:0] _T_660; // @[Lookup.scala 11:37:@1282.4]
  wire [2:0] _T_661; // @[Lookup.scala 11:37:@1283.4]
  wire [2:0] _T_662; // @[Lookup.scala 11:37:@1284.4]
  wire [2:0] _T_663; // @[Lookup.scala 11:37:@1285.4]
  wire [2:0] ctlsig_6; // @[Lookup.scala 11:37:@1286.4]
  wire [1:0] _T_664; // @[Lookup.scala 11:37:@1287.4]
  wire [1:0] _T_665; // @[Lookup.scala 11:37:@1288.4]
  wire [1:0] _T_666; // @[Lookup.scala 11:37:@1289.4]
  wire [1:0] _T_667; // @[Lookup.scala 11:37:@1290.4]
  wire [1:0] _T_668; // @[Lookup.scala 11:37:@1291.4]
  wire [1:0] _T_669; // @[Lookup.scala 11:37:@1292.4]
  wire [1:0] _T_670; // @[Lookup.scala 11:37:@1293.4]
  wire [1:0] _T_671; // @[Lookup.scala 11:37:@1294.4]
  wire [1:0] _T_672; // @[Lookup.scala 11:37:@1295.4]
  wire [1:0] _T_673; // @[Lookup.scala 11:37:@1296.4]
  wire [1:0] _T_674; // @[Lookup.scala 11:37:@1297.4]
  wire [1:0] _T_675; // @[Lookup.scala 11:37:@1298.4]
  wire [1:0] _T_676; // @[Lookup.scala 11:37:@1299.4]
  wire [1:0] _T_677; // @[Lookup.scala 11:37:@1300.4]
  wire [1:0] _T_678; // @[Lookup.scala 11:37:@1301.4]
  wire [1:0] _T_679; // @[Lookup.scala 11:37:@1302.4]
  wire [1:0] _T_680; // @[Lookup.scala 11:37:@1303.4]
  wire [1:0] _T_681; // @[Lookup.scala 11:37:@1304.4]
  wire [1:0] _T_682; // @[Lookup.scala 11:37:@1305.4]
  wire [1:0] _T_683; // @[Lookup.scala 11:37:@1306.4]
  wire [1:0] _T_684; // @[Lookup.scala 11:37:@1307.4]
  wire [1:0] _T_685; // @[Lookup.scala 11:37:@1308.4]
  wire [1:0] _T_686; // @[Lookup.scala 11:37:@1309.4]
  wire [1:0] _T_687; // @[Lookup.scala 11:37:@1310.4]
  wire [1:0] _T_688; // @[Lookup.scala 11:37:@1311.4]
  wire [1:0] _T_689; // @[Lookup.scala 11:37:@1312.4]
  wire [1:0] _T_690; // @[Lookup.scala 11:37:@1313.4]
  wire [1:0] _T_691; // @[Lookup.scala 11:37:@1314.4]
  wire [1:0] _T_692; // @[Lookup.scala 11:37:@1315.4]
  wire [1:0] _T_693; // @[Lookup.scala 11:37:@1316.4]
  wire [1:0] _T_694; // @[Lookup.scala 11:37:@1317.4]
  wire [1:0] _T_695; // @[Lookup.scala 11:37:@1318.4]
  wire [1:0] _T_696; // @[Lookup.scala 11:37:@1319.4]
  wire [1:0] _T_697; // @[Lookup.scala 11:37:@1320.4]
  wire [1:0] _T_698; // @[Lookup.scala 11:37:@1321.4]
  wire [1:0] _T_699; // @[Lookup.scala 11:37:@1322.4]
  wire [1:0] _T_700; // @[Lookup.scala 11:37:@1323.4]
  wire [1:0] _T_701; // @[Lookup.scala 11:37:@1324.4]
  wire [1:0] _T_702; // @[Lookup.scala 11:37:@1325.4]
  wire [1:0] _T_703; // @[Lookup.scala 11:37:@1326.4]
  wire [1:0] _T_704; // @[Lookup.scala 11:37:@1327.4]
  wire [1:0] _T_705; // @[Lookup.scala 11:37:@1328.4]
  wire [1:0] _T_706; // @[Lookup.scala 11:37:@1329.4]
  wire [1:0] _T_707; // @[Lookup.scala 11:37:@1330.4]
  wire [1:0] _T_708; // @[Lookup.scala 11:37:@1331.4]
  wire [1:0] _T_709; // @[Lookup.scala 11:37:@1332.4]
  wire [1:0] _T_710; // @[Lookup.scala 11:37:@1333.4]
  wire [1:0] _T_711; // @[Lookup.scala 11:37:@1334.4]
  wire [1:0] _T_712; // @[Lookup.scala 11:37:@1335.4]
  wire [1:0] ctlsig_7; // @[Lookup.scala 11:37:@1336.4]
  wire [2:0] _T_753; // @[Lookup.scala 11:37:@1377.4]
  wire [2:0] _T_754; // @[Lookup.scala 11:37:@1378.4]
  wire [2:0] _T_755; // @[Lookup.scala 11:37:@1379.4]
  wire [2:0] _T_756; // @[Lookup.scala 11:37:@1380.4]
  wire [2:0] _T_757; // @[Lookup.scala 11:37:@1381.4]
  wire [2:0] _T_758; // @[Lookup.scala 11:37:@1382.4]
  wire [2:0] _T_759; // @[Lookup.scala 11:37:@1383.4]
  wire [2:0] _T_760; // @[Lookup.scala 11:37:@1384.4]
  wire [2:0] _T_761; // @[Lookup.scala 11:37:@1385.4]
  wire [2:0] br_sel; // @[Lookup.scala 11:37:@1386.4]
  wire [1:0] _T_769; // @[Lookup.scala 11:37:@1394.4]
  wire [1:0] _T_770; // @[Lookup.scala 11:37:@1395.4]
  wire [1:0] _T_771; // @[Lookup.scala 11:37:@1396.4]
  wire [1:0] _T_772; // @[Lookup.scala 11:37:@1397.4]
  wire [1:0] _T_773; // @[Lookup.scala 11:37:@1398.4]
  wire [1:0] _T_774; // @[Lookup.scala 11:37:@1399.4]
  wire [1:0] _T_775; // @[Lookup.scala 11:37:@1400.4]
  wire [1:0] _T_776; // @[Lookup.scala 11:37:@1401.4]
  wire [1:0] _T_777; // @[Lookup.scala 11:37:@1402.4]
  wire [1:0] _T_778; // @[Lookup.scala 11:37:@1403.4]
  wire [1:0] _T_779; // @[Lookup.scala 11:37:@1404.4]
  wire [1:0] _T_780; // @[Lookup.scala 11:37:@1405.4]
  wire [1:0] _T_781; // @[Lookup.scala 11:37:@1406.4]
  wire [1:0] _T_782; // @[Lookup.scala 11:37:@1407.4]
  wire [1:0] _T_783; // @[Lookup.scala 11:37:@1408.4]
  wire [1:0] _T_784; // @[Lookup.scala 11:37:@1409.4]
  wire [1:0] _T_785; // @[Lookup.scala 11:37:@1410.4]
  wire [1:0] _T_786; // @[Lookup.scala 11:37:@1411.4]
  wire [1:0] _T_787; // @[Lookup.scala 11:37:@1412.4]
  wire [1:0] _T_788; // @[Lookup.scala 11:37:@1413.4]
  wire [1:0] _T_789; // @[Lookup.scala 11:37:@1414.4]
  wire [1:0] _T_790; // @[Lookup.scala 11:37:@1415.4]
  wire [1:0] _T_791; // @[Lookup.scala 11:37:@1416.4]
  wire [1:0] _T_792; // @[Lookup.scala 11:37:@1417.4]
  wire [1:0] _T_793; // @[Lookup.scala 11:37:@1418.4]
  wire [1:0] _T_794; // @[Lookup.scala 11:37:@1419.4]
  wire [1:0] _T_795; // @[Lookup.scala 11:37:@1420.4]
  wire [1:0] _T_796; // @[Lookup.scala 11:37:@1421.4]
  wire [1:0] _T_797; // @[Lookup.scala 11:37:@1422.4]
  wire [1:0] _T_798; // @[Lookup.scala 11:37:@1423.4]
  wire [1:0] _T_799; // @[Lookup.scala 11:37:@1424.4]
  wire [1:0] _T_800; // @[Lookup.scala 11:37:@1425.4]
  wire [1:0] _T_801; // @[Lookup.scala 11:37:@1426.4]
  wire [1:0] _T_802; // @[Lookup.scala 11:37:@1427.4]
  wire [1:0] _T_803; // @[Lookup.scala 11:37:@1428.4]
  wire [1:0] _T_804; // @[Lookup.scala 11:37:@1429.4]
  wire [1:0] _T_805; // @[Lookup.scala 11:37:@1430.4]
  wire [1:0] _T_806; // @[Lookup.scala 11:37:@1431.4]
  wire [1:0] _T_807; // @[Lookup.scala 11:37:@1432.4]
  wire [1:0] _T_808; // @[Lookup.scala 11:37:@1433.4]
  wire [1:0] _T_809; // @[Lookup.scala 11:37:@1434.4]
  wire [1:0] _T_810; // @[Lookup.scala 11:37:@1435.4]
  wire [1:0] ctlsig_9; // @[Lookup.scala 11:37:@1436.4]
  wire [2:0] _T_811; // @[Lookup.scala 11:37:@1437.4]
  wire [2:0] _T_812; // @[Lookup.scala 11:37:@1438.4]
  wire [2:0] _T_813; // @[Lookup.scala 11:37:@1439.4]
  wire [2:0] _T_814; // @[Lookup.scala 11:37:@1440.4]
  wire [2:0] _T_815; // @[Lookup.scala 11:37:@1441.4]
  wire [2:0] _T_816; // @[Lookup.scala 11:37:@1442.4]
  wire [2:0] _T_817; // @[Lookup.scala 11:37:@1443.4]
  wire [2:0] _T_818; // @[Lookup.scala 11:37:@1444.4]
  wire [2:0] _T_819; // @[Lookup.scala 11:37:@1445.4]
  wire [2:0] _T_820; // @[Lookup.scala 11:37:@1446.4]
  wire [2:0] _T_821; // @[Lookup.scala 11:37:@1447.4]
  wire [2:0] _T_822; // @[Lookup.scala 11:37:@1448.4]
  wire [2:0] _T_823; // @[Lookup.scala 11:37:@1449.4]
  wire [2:0] _T_824; // @[Lookup.scala 11:37:@1450.4]
  wire [2:0] _T_825; // @[Lookup.scala 11:37:@1451.4]
  wire [2:0] _T_826; // @[Lookup.scala 11:37:@1452.4]
  wire [2:0] _T_827; // @[Lookup.scala 11:37:@1453.4]
  wire [2:0] _T_828; // @[Lookup.scala 11:37:@1454.4]
  wire [2:0] _T_829; // @[Lookup.scala 11:37:@1455.4]
  wire [2:0] _T_830; // @[Lookup.scala 11:37:@1456.4]
  wire [2:0] _T_831; // @[Lookup.scala 11:37:@1457.4]
  wire [2:0] _T_832; // @[Lookup.scala 11:37:@1458.4]
  wire [2:0] _T_833; // @[Lookup.scala 11:37:@1459.4]
  wire [2:0] _T_834; // @[Lookup.scala 11:37:@1460.4]
  wire [2:0] _T_835; // @[Lookup.scala 11:37:@1461.4]
  wire [2:0] _T_836; // @[Lookup.scala 11:37:@1462.4]
  wire [2:0] _T_837; // @[Lookup.scala 11:37:@1463.4]
  wire [2:0] _T_838; // @[Lookup.scala 11:37:@1464.4]
  wire [2:0] _T_839; // @[Lookup.scala 11:37:@1465.4]
  wire [2:0] _T_840; // @[Lookup.scala 11:37:@1466.4]
  wire [2:0] _T_841; // @[Lookup.scala 11:37:@1467.4]
  wire [2:0] _T_842; // @[Lookup.scala 11:37:@1468.4]
  wire [2:0] _T_843; // @[Lookup.scala 11:37:@1469.4]
  wire [2:0] _T_844; // @[Lookup.scala 11:37:@1470.4]
  wire [2:0] _T_845; // @[Lookup.scala 11:37:@1471.4]
  wire [2:0] _T_846; // @[Lookup.scala 11:37:@1472.4]
  wire [2:0] _T_847; // @[Lookup.scala 11:37:@1473.4]
  wire [2:0] _T_848; // @[Lookup.scala 11:37:@1474.4]
  wire [2:0] _T_849; // @[Lookup.scala 11:37:@1475.4]
  wire [2:0] _T_850; // @[Lookup.scala 11:37:@1476.4]
  wire [2:0] _T_851; // @[Lookup.scala 11:37:@1477.4]
  wire [2:0] _T_852; // @[Lookup.scala 11:37:@1478.4]
  wire [2:0] _T_853; // @[Lookup.scala 11:37:@1479.4]
  wire [2:0] _T_854; // @[Lookup.scala 11:37:@1480.4]
  wire [2:0] _T_855; // @[Lookup.scala 11:37:@1481.4]
  wire [2:0] _T_856; // @[Lookup.scala 11:37:@1482.4]
  wire [2:0] _T_857; // @[Lookup.scala 11:37:@1483.4]
  wire [2:0] _T_858; // @[Lookup.scala 11:37:@1484.4]
  wire [2:0] _T_859; // @[Lookup.scala 11:37:@1485.4]
  wire [2:0] csr_cmd; // @[Lookup.scala 11:37:@1486.4]
  wire  _T_861; // @[Lookup.scala 11:37:@1488.4]
  wire  _T_862; // @[Lookup.scala 11:37:@1489.4]
  wire  _T_863; // @[Lookup.scala 11:37:@1490.4]
  wire  _T_864; // @[Lookup.scala 11:37:@1491.4]
  wire  _T_865; // @[Lookup.scala 11:37:@1492.4]
  wire  _T_866; // @[Lookup.scala 11:37:@1493.4]
  wire  _T_867; // @[Lookup.scala 11:37:@1494.4]
  wire  _T_868; // @[Lookup.scala 11:37:@1495.4]
  wire  _T_869; // @[Lookup.scala 11:37:@1496.4]
  wire  _T_870; // @[Lookup.scala 11:37:@1497.4]
  wire  _T_871; // @[Lookup.scala 11:37:@1498.4]
  wire  _T_872; // @[Lookup.scala 11:37:@1499.4]
  wire  _T_873; // @[Lookup.scala 11:37:@1500.4]
  wire  _T_874; // @[Lookup.scala 11:37:@1501.4]
  wire  _T_875; // @[Lookup.scala 11:37:@1502.4]
  wire  _T_876; // @[Lookup.scala 11:37:@1503.4]
  wire  _T_877; // @[Lookup.scala 11:37:@1504.4]
  wire  _T_878; // @[Lookup.scala 11:37:@1505.4]
  wire  _T_879; // @[Lookup.scala 11:37:@1506.4]
  wire  _T_880; // @[Lookup.scala 11:37:@1507.4]
  wire  _T_881; // @[Lookup.scala 11:37:@1508.4]
  wire  _T_882; // @[Lookup.scala 11:37:@1509.4]
  wire  _T_883; // @[Lookup.scala 11:37:@1510.4]
  wire  _T_884; // @[Lookup.scala 11:37:@1511.4]
  wire  _T_885; // @[Lookup.scala 11:37:@1512.4]
  wire  _T_886; // @[Lookup.scala 11:37:@1513.4]
  wire  _T_887; // @[Lookup.scala 11:37:@1514.4]
  wire  _T_888; // @[Lookup.scala 11:37:@1515.4]
  wire  _T_889; // @[Lookup.scala 11:37:@1516.4]
  wire  _T_890; // @[Lookup.scala 11:37:@1517.4]
  wire  _T_891; // @[Lookup.scala 11:37:@1518.4]
  wire  _T_892; // @[Lookup.scala 11:37:@1519.4]
  wire  _T_893; // @[Lookup.scala 11:37:@1520.4]
  wire  _T_894; // @[Lookup.scala 11:37:@1521.4]
  wire  _T_895; // @[Lookup.scala 11:37:@1522.4]
  wire  _T_896; // @[Lookup.scala 11:37:@1523.4]
  wire  _T_897; // @[Lookup.scala 11:37:@1524.4]
  wire  _T_898; // @[Lookup.scala 11:37:@1525.4]
  wire  _T_899; // @[Lookup.scala 11:37:@1526.4]
  wire  _T_900; // @[Lookup.scala 11:37:@1527.4]
  wire  _T_901; // @[Lookup.scala 11:37:@1528.4]
  wire  _T_902; // @[Lookup.scala 11:37:@1529.4]
  wire  _T_903; // @[Lookup.scala 11:37:@1530.4]
  wire  _T_904; // @[Lookup.scala 11:37:@1531.4]
  wire  _T_905; // @[Lookup.scala 11:37:@1532.4]
  wire  _T_906; // @[Lookup.scala 11:37:@1533.4]
  wire  _T_907; // @[Lookup.scala 11:37:@1534.4]
  wire  _T_908; // @[Lookup.scala 11:37:@1535.4]
  wire  ctlsig_11; // @[Lookup.scala 11:37:@1536.4]
  wire  _T_909; // @[rvcpath.scala 134:39:@1544.4]
  wire [1:0] _T_910; // @[rvcpath.scala 134:25:@1545.4]
  wire  _T_911; // @[rvcpath.scala 139:33:@1550.4]
  wire [3:0] _T_913; // @[rvcpath.scala 140:25:@1552.4]
  assign _T_123 = io_d2c_inst & 32'h7f; // @[Lookup.scala 9:38:@837.4]
  assign _T_124 = 32'h37 == _T_123; // @[Lookup.scala 9:38:@838.4]
  assign _T_128 = 32'h17 == _T_123; // @[Lookup.scala 9:38:@840.4]
  assign _T_132 = 32'h6f == _T_123; // @[Lookup.scala 9:38:@842.4]
  assign _T_135 = io_d2c_inst & 32'h707f; // @[Lookup.scala 9:38:@843.4]
  assign _T_136 = 32'h67 == _T_135; // @[Lookup.scala 9:38:@844.4]
  assign _T_140 = 32'h63 == _T_135; // @[Lookup.scala 9:38:@846.4]
  assign _T_144 = 32'h1063 == _T_135; // @[Lookup.scala 9:38:@848.4]
  assign _T_148 = 32'h4063 == _T_135; // @[Lookup.scala 9:38:@850.4]
  assign _T_152 = 32'h5063 == _T_135; // @[Lookup.scala 9:38:@852.4]
  assign _T_156 = 32'h6063 == _T_135; // @[Lookup.scala 9:38:@854.4]
  assign _T_160 = 32'h7063 == _T_135; // @[Lookup.scala 9:38:@856.4]
  assign _T_164 = 32'h3 == _T_135; // @[Lookup.scala 9:38:@858.4]
  assign _T_168 = 32'h1003 == _T_135; // @[Lookup.scala 9:38:@860.4]
  assign _T_172 = 32'h2003 == _T_135; // @[Lookup.scala 9:38:@862.4]
  assign _T_176 = 32'h4003 == _T_135; // @[Lookup.scala 9:38:@864.4]
  assign _T_180 = 32'h5003 == _T_135; // @[Lookup.scala 9:38:@866.4]
  assign _T_184 = 32'h23 == _T_135; // @[Lookup.scala 9:38:@868.4]
  assign _T_188 = 32'h1023 == _T_135; // @[Lookup.scala 9:38:@870.4]
  assign _T_192 = 32'h2023 == _T_135; // @[Lookup.scala 9:38:@872.4]
  assign _T_196 = 32'h13 == _T_135; // @[Lookup.scala 9:38:@874.4]
  assign _T_200 = 32'h2013 == _T_135; // @[Lookup.scala 9:38:@876.4]
  assign _T_204 = 32'h3013 == _T_135; // @[Lookup.scala 9:38:@878.4]
  assign _T_208 = 32'h4013 == _T_135; // @[Lookup.scala 9:38:@880.4]
  assign _T_212 = 32'h6013 == _T_135; // @[Lookup.scala 9:38:@882.4]
  assign _T_216 = 32'h7013 == _T_135; // @[Lookup.scala 9:38:@884.4]
  assign _T_219 = io_d2c_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@885.4]
  assign _T_220 = 32'h1013 == _T_219; // @[Lookup.scala 9:38:@886.4]
  assign _T_224 = 32'h5013 == _T_219; // @[Lookup.scala 9:38:@888.4]
  assign _T_228 = 32'h40005013 == _T_219; // @[Lookup.scala 9:38:@890.4]
  assign _T_232 = 32'h33 == _T_219; // @[Lookup.scala 9:38:@892.4]
  assign _T_236 = 32'h40000033 == _T_219; // @[Lookup.scala 9:38:@894.4]
  assign _T_240 = 32'h1033 == _T_219; // @[Lookup.scala 9:38:@896.4]
  assign _T_244 = 32'h2033 == _T_219; // @[Lookup.scala 9:38:@898.4]
  assign _T_248 = 32'h3033 == _T_219; // @[Lookup.scala 9:38:@900.4]
  assign _T_252 = 32'h4033 == _T_219; // @[Lookup.scala 9:38:@902.4]
  assign _T_256 = 32'h5033 == _T_219; // @[Lookup.scala 9:38:@904.4]
  assign _T_260 = 32'h40005033 == _T_219; // @[Lookup.scala 9:38:@906.4]
  assign _T_264 = 32'h6033 == _T_219; // @[Lookup.scala 9:38:@908.4]
  assign _T_268 = 32'h7033 == _T_219; // @[Lookup.scala 9:38:@910.4]
  assign _T_272 = 32'h1073 == _T_135; // @[Lookup.scala 9:38:@912.4]
  assign _T_276 = 32'h2073 == _T_135; // @[Lookup.scala 9:38:@914.4]
  assign _T_280 = 32'h3073 == _T_135; // @[Lookup.scala 9:38:@916.4]
  assign _T_284 = 32'h5073 == _T_135; // @[Lookup.scala 9:38:@918.4]
  assign _T_288 = 32'h6073 == _T_135; // @[Lookup.scala 9:38:@920.4]
  assign _T_292 = 32'h7073 == _T_135; // @[Lookup.scala 9:38:@922.4]
  assign _T_295 = io_d2c_inst & 32'hf00fffff; // @[Lookup.scala 9:38:@923.4]
  assign _T_296 = 32'hf == _T_295; // @[Lookup.scala 9:38:@924.4]
  assign _T_300 = 32'h100f == io_d2c_inst; // @[Lookup.scala 9:38:@926.4]
  assign _T_304 = 32'h73 == io_d2c_inst; // @[Lookup.scala 9:38:@928.4]
  assign _T_308 = 32'h100073 == io_d2c_inst; // @[Lookup.scala 9:38:@930.4]
  assign _T_312 = 32'h30200073 == io_d2c_inst; // @[Lookup.scala 9:38:@932.4]
  assign _T_316 = 32'h10500073 == io_d2c_inst; // @[Lookup.scala 9:38:@934.4]
  assign _T_320 = 32'h7b200073 == io_d2c_inst; // @[Lookup.scala 9:38:@936.4]
  assign _T_334 = _T_268 ? 4'h7 : 4'hf; // @[Lookup.scala 11:37:@950.4]
  assign _T_335 = _T_264 ? 4'h6 : _T_334; // @[Lookup.scala 11:37:@951.4]
  assign _T_336 = _T_260 ? 4'hd : _T_335; // @[Lookup.scala 11:37:@952.4]
  assign _T_337 = _T_256 ? 4'h5 : _T_336; // @[Lookup.scala 11:37:@953.4]
  assign _T_338 = _T_252 ? 4'h4 : _T_337; // @[Lookup.scala 11:37:@954.4]
  assign _T_339 = _T_248 ? 4'h3 : _T_338; // @[Lookup.scala 11:37:@955.4]
  assign _T_340 = _T_244 ? 4'h2 : _T_339; // @[Lookup.scala 11:37:@956.4]
  assign _T_341 = _T_240 ? 4'h1 : _T_340; // @[Lookup.scala 11:37:@957.4]
  assign _T_342 = _T_236 ? 4'h8 : _T_341; // @[Lookup.scala 11:37:@958.4]
  assign _T_343 = _T_232 ? 4'h0 : _T_342; // @[Lookup.scala 11:37:@959.4]
  assign _T_344 = _T_228 ? 4'hd : _T_343; // @[Lookup.scala 11:37:@960.4]
  assign _T_345 = _T_224 ? 4'h5 : _T_344; // @[Lookup.scala 11:37:@961.4]
  assign _T_346 = _T_220 ? 4'h1 : _T_345; // @[Lookup.scala 11:37:@962.4]
  assign _T_347 = _T_216 ? 4'h7 : _T_346; // @[Lookup.scala 11:37:@963.4]
  assign _T_348 = _T_212 ? 4'h6 : _T_347; // @[Lookup.scala 11:37:@964.4]
  assign _T_349 = _T_208 ? 4'h4 : _T_348; // @[Lookup.scala 11:37:@965.4]
  assign _T_350 = _T_204 ? 4'h3 : _T_349; // @[Lookup.scala 11:37:@966.4]
  assign _T_351 = _T_200 ? 4'h2 : _T_350; // @[Lookup.scala 11:37:@967.4]
  assign _T_352 = _T_196 ? 4'h0 : _T_351; // @[Lookup.scala 11:37:@968.4]
  assign _T_353 = _T_192 ? 4'h0 : _T_352; // @[Lookup.scala 11:37:@969.4]
  assign _T_354 = _T_188 ? 4'h0 : _T_353; // @[Lookup.scala 11:37:@970.4]
  assign _T_355 = _T_184 ? 4'h0 : _T_354; // @[Lookup.scala 11:37:@971.4]
  assign _T_356 = _T_180 ? 4'h0 : _T_355; // @[Lookup.scala 11:37:@972.4]
  assign _T_357 = _T_176 ? 4'h0 : _T_356; // @[Lookup.scala 11:37:@973.4]
  assign _T_358 = _T_172 ? 4'h0 : _T_357; // @[Lookup.scala 11:37:@974.4]
  assign _T_359 = _T_168 ? 4'h0 : _T_358; // @[Lookup.scala 11:37:@975.4]
  assign _T_360 = _T_164 ? 4'h0 : _T_359; // @[Lookup.scala 11:37:@976.4]
  assign _T_361 = _T_160 ? 4'h0 : _T_360; // @[Lookup.scala 11:37:@977.4]
  assign _T_362 = _T_156 ? 4'h0 : _T_361; // @[Lookup.scala 11:37:@978.4]
  assign _T_363 = _T_152 ? 4'h0 : _T_362; // @[Lookup.scala 11:37:@979.4]
  assign _T_364 = _T_148 ? 4'h0 : _T_363; // @[Lookup.scala 11:37:@980.4]
  assign _T_365 = _T_144 ? 4'h0 : _T_364; // @[Lookup.scala 11:37:@981.4]
  assign _T_366 = _T_140 ? 4'h0 : _T_365; // @[Lookup.scala 11:37:@982.4]
  assign _T_367 = _T_136 ? 4'h0 : _T_366; // @[Lookup.scala 11:37:@983.4]
  assign _T_368 = _T_132 ? 4'h0 : _T_367; // @[Lookup.scala 11:37:@984.4]
  assign _T_369 = _T_128 ? 4'h0 : _T_368; // @[Lookup.scala 11:37:@985.4]
  assign alu_func = _T_124 ? 4'hb : _T_369; // @[Lookup.scala 11:37:@986.4]
  assign _T_383 = _T_268 ? 3'h0 : 3'h7; // @[Lookup.scala 11:37:@1000.4]
  assign _T_384 = _T_264 ? 3'h0 : _T_383; // @[Lookup.scala 11:37:@1001.4]
  assign _T_385 = _T_260 ? 3'h0 : _T_384; // @[Lookup.scala 11:37:@1002.4]
  assign _T_386 = _T_256 ? 3'h0 : _T_385; // @[Lookup.scala 11:37:@1003.4]
  assign _T_387 = _T_252 ? 3'h0 : _T_386; // @[Lookup.scala 11:37:@1004.4]
  assign _T_388 = _T_248 ? 3'h0 : _T_387; // @[Lookup.scala 11:37:@1005.4]
  assign _T_389 = _T_244 ? 3'h0 : _T_388; // @[Lookup.scala 11:37:@1006.4]
  assign _T_390 = _T_240 ? 3'h0 : _T_389; // @[Lookup.scala 11:37:@1007.4]
  assign _T_391 = _T_236 ? 3'h0 : _T_390; // @[Lookup.scala 11:37:@1008.4]
  assign _T_392 = _T_232 ? 3'h0 : _T_391; // @[Lookup.scala 11:37:@1009.4]
  assign _T_393 = _T_228 ? 3'h1 : _T_392; // @[Lookup.scala 11:37:@1010.4]
  assign _T_394 = _T_224 ? 3'h1 : _T_393; // @[Lookup.scala 11:37:@1011.4]
  assign _T_395 = _T_220 ? 3'h1 : _T_394; // @[Lookup.scala 11:37:@1012.4]
  assign _T_396 = _T_216 ? 3'h1 : _T_395; // @[Lookup.scala 11:37:@1013.4]
  assign _T_397 = _T_212 ? 3'h1 : _T_396; // @[Lookup.scala 11:37:@1014.4]
  assign _T_398 = _T_208 ? 3'h1 : _T_397; // @[Lookup.scala 11:37:@1015.4]
  assign _T_399 = _T_204 ? 3'h1 : _T_398; // @[Lookup.scala 11:37:@1016.4]
  assign _T_400 = _T_200 ? 3'h1 : _T_399; // @[Lookup.scala 11:37:@1017.4]
  assign _T_401 = _T_196 ? 3'h1 : _T_400; // @[Lookup.scala 11:37:@1018.4]
  assign _T_402 = _T_192 ? 3'h2 : _T_401; // @[Lookup.scala 11:37:@1019.4]
  assign _T_403 = _T_188 ? 3'h2 : _T_402; // @[Lookup.scala 11:37:@1020.4]
  assign _T_404 = _T_184 ? 3'h2 : _T_403; // @[Lookup.scala 11:37:@1021.4]
  assign _T_405 = _T_180 ? 3'h1 : _T_404; // @[Lookup.scala 11:37:@1022.4]
  assign _T_406 = _T_176 ? 3'h1 : _T_405; // @[Lookup.scala 11:37:@1023.4]
  assign _T_407 = _T_172 ? 3'h1 : _T_406; // @[Lookup.scala 11:37:@1024.4]
  assign _T_408 = _T_168 ? 3'h1 : _T_407; // @[Lookup.scala 11:37:@1025.4]
  assign _T_409 = _T_164 ? 3'h1 : _T_408; // @[Lookup.scala 11:37:@1026.4]
  assign _T_410 = _T_160 ? 3'h3 : _T_409; // @[Lookup.scala 11:37:@1027.4]
  assign _T_411 = _T_156 ? 3'h3 : _T_410; // @[Lookup.scala 11:37:@1028.4]
  assign _T_412 = _T_152 ? 3'h3 : _T_411; // @[Lookup.scala 11:37:@1029.4]
  assign _T_413 = _T_148 ? 3'h3 : _T_412; // @[Lookup.scala 11:37:@1030.4]
  assign _T_414 = _T_144 ? 3'h3 : _T_413; // @[Lookup.scala 11:37:@1031.4]
  assign _T_415 = _T_140 ? 3'h3 : _T_414; // @[Lookup.scala 11:37:@1032.4]
  assign _T_416 = _T_136 ? 3'h1 : _T_415; // @[Lookup.scala 11:37:@1033.4]
  assign _T_417 = _T_132 ? 3'h5 : _T_416; // @[Lookup.scala 11:37:@1034.4]
  assign _T_418 = _T_128 ? 3'h4 : _T_417; // @[Lookup.scala 11:37:@1035.4]
  assign ctlsig_1 = _T_124 ? 3'h4 : _T_418; // @[Lookup.scala 11:37:@1036.4]
  assign _T_427 = _T_288 ? 1'h1 : _T_292; // @[Lookup.scala 11:37:@1045.4]
  assign _T_428 = _T_284 ? 1'h1 : _T_427; // @[Lookup.scala 11:37:@1046.4]
  assign _T_429 = _T_280 ? 1'h1 : _T_428; // @[Lookup.scala 11:37:@1047.4]
  assign _T_430 = _T_276 ? 1'h1 : _T_429; // @[Lookup.scala 11:37:@1048.4]
  assign _T_431 = _T_272 ? 1'h1 : _T_430; // @[Lookup.scala 11:37:@1049.4]
  assign _T_432 = _T_268 ? 1'h1 : _T_431; // @[Lookup.scala 11:37:@1050.4]
  assign _T_433 = _T_264 ? 1'h1 : _T_432; // @[Lookup.scala 11:37:@1051.4]
  assign _T_434 = _T_260 ? 1'h1 : _T_433; // @[Lookup.scala 11:37:@1052.4]
  assign _T_435 = _T_256 ? 1'h1 : _T_434; // @[Lookup.scala 11:37:@1053.4]
  assign _T_436 = _T_252 ? 1'h1 : _T_435; // @[Lookup.scala 11:37:@1054.4]
  assign _T_437 = _T_248 ? 1'h1 : _T_436; // @[Lookup.scala 11:37:@1055.4]
  assign _T_438 = _T_244 ? 1'h1 : _T_437; // @[Lookup.scala 11:37:@1056.4]
  assign _T_439 = _T_240 ? 1'h1 : _T_438; // @[Lookup.scala 11:37:@1057.4]
  assign _T_440 = _T_236 ? 1'h1 : _T_439; // @[Lookup.scala 11:37:@1058.4]
  assign _T_441 = _T_232 ? 1'h1 : _T_440; // @[Lookup.scala 11:37:@1059.4]
  assign _T_442 = _T_228 ? 1'h1 : _T_441; // @[Lookup.scala 11:37:@1060.4]
  assign _T_443 = _T_224 ? 1'h1 : _T_442; // @[Lookup.scala 11:37:@1061.4]
  assign _T_444 = _T_220 ? 1'h1 : _T_443; // @[Lookup.scala 11:37:@1062.4]
  assign _T_445 = _T_216 ? 1'h1 : _T_444; // @[Lookup.scala 11:37:@1063.4]
  assign _T_446 = _T_212 ? 1'h1 : _T_445; // @[Lookup.scala 11:37:@1064.4]
  assign _T_447 = _T_208 ? 1'h1 : _T_446; // @[Lookup.scala 11:37:@1065.4]
  assign _T_448 = _T_204 ? 1'h1 : _T_447; // @[Lookup.scala 11:37:@1066.4]
  assign _T_449 = _T_200 ? 1'h1 : _T_448; // @[Lookup.scala 11:37:@1067.4]
  assign _T_450 = _T_196 ? 1'h1 : _T_449; // @[Lookup.scala 11:37:@1068.4]
  assign _T_451 = _T_192 ? 1'h0 : _T_450; // @[Lookup.scala 11:37:@1069.4]
  assign _T_452 = _T_188 ? 1'h0 : _T_451; // @[Lookup.scala 11:37:@1070.4]
  assign _T_453 = _T_184 ? 1'h0 : _T_452; // @[Lookup.scala 11:37:@1071.4]
  assign _T_454 = _T_180 ? 1'h1 : _T_453; // @[Lookup.scala 11:37:@1072.4]
  assign _T_455 = _T_176 ? 1'h1 : _T_454; // @[Lookup.scala 11:37:@1073.4]
  assign _T_456 = _T_172 ? 1'h1 : _T_455; // @[Lookup.scala 11:37:@1074.4]
  assign _T_457 = _T_168 ? 1'h1 : _T_456; // @[Lookup.scala 11:37:@1075.4]
  assign _T_458 = _T_164 ? 1'h1 : _T_457; // @[Lookup.scala 11:37:@1076.4]
  assign _T_459 = _T_160 ? 1'h0 : _T_458; // @[Lookup.scala 11:37:@1077.4]
  assign _T_460 = _T_156 ? 1'h0 : _T_459; // @[Lookup.scala 11:37:@1078.4]
  assign _T_461 = _T_152 ? 1'h0 : _T_460; // @[Lookup.scala 11:37:@1079.4]
  assign _T_462 = _T_148 ? 1'h0 : _T_461; // @[Lookup.scala 11:37:@1080.4]
  assign _T_463 = _T_144 ? 1'h0 : _T_462; // @[Lookup.scala 11:37:@1081.4]
  assign _T_464 = _T_140 ? 1'h0 : _T_463; // @[Lookup.scala 11:37:@1082.4]
  assign _T_465 = _T_136 ? 1'h1 : _T_464; // @[Lookup.scala 11:37:@1083.4]
  assign _T_466 = _T_132 ? 1'h1 : _T_465; // @[Lookup.scala 11:37:@1084.4]
  assign _T_467 = _T_128 ? 1'h1 : _T_466; // @[Lookup.scala 11:37:@1085.4]
  assign ctlsig_2 = _T_124 ? 1'h1 : _T_467; // @[Lookup.scala 11:37:@1086.4]
  assign _T_501 = _T_188 ? 1'h1 : _T_192; // @[Lookup.scala 11:37:@1120.4]
  assign _T_502 = _T_184 ? 1'h1 : _T_501; // @[Lookup.scala 11:37:@1121.4]
  assign _T_503 = _T_180 ? 1'h0 : _T_502; // @[Lookup.scala 11:37:@1122.4]
  assign _T_504 = _T_176 ? 1'h0 : _T_503; // @[Lookup.scala 11:37:@1123.4]
  assign _T_505 = _T_172 ? 1'h0 : _T_504; // @[Lookup.scala 11:37:@1124.4]
  assign _T_506 = _T_168 ? 1'h0 : _T_505; // @[Lookup.scala 11:37:@1125.4]
  assign _T_507 = _T_164 ? 1'h0 : _T_506; // @[Lookup.scala 11:37:@1126.4]
  assign _T_508 = _T_160 ? 1'h0 : _T_507; // @[Lookup.scala 11:37:@1127.4]
  assign _T_509 = _T_156 ? 1'h0 : _T_508; // @[Lookup.scala 11:37:@1128.4]
  assign _T_510 = _T_152 ? 1'h0 : _T_509; // @[Lookup.scala 11:37:@1129.4]
  assign _T_511 = _T_148 ? 1'h0 : _T_510; // @[Lookup.scala 11:37:@1130.4]
  assign _T_512 = _T_144 ? 1'h0 : _T_511; // @[Lookup.scala 11:37:@1131.4]
  assign _T_513 = _T_140 ? 1'h0 : _T_512; // @[Lookup.scala 11:37:@1132.4]
  assign _T_514 = _T_136 ? 1'h0 : _T_513; // @[Lookup.scala 11:37:@1133.4]
  assign _T_515 = _T_132 ? 1'h0 : _T_514; // @[Lookup.scala 11:37:@1134.4]
  assign _T_516 = _T_128 ? 1'h0 : _T_515; // @[Lookup.scala 11:37:@1135.4]
  assign ctlsig_3 = _T_124 ? 1'h0 : _T_516; // @[Lookup.scala 11:37:@1136.4]
  assign _T_552 = _T_180 ? 1'h1 : _T_502; // @[Lookup.scala 11:37:@1172.4]
  assign _T_553 = _T_176 ? 1'h1 : _T_552; // @[Lookup.scala 11:37:@1173.4]
  assign _T_554 = _T_172 ? 1'h1 : _T_553; // @[Lookup.scala 11:37:@1174.4]
  assign _T_555 = _T_168 ? 1'h1 : _T_554; // @[Lookup.scala 11:37:@1175.4]
  assign _T_556 = _T_164 ? 1'h1 : _T_555; // @[Lookup.scala 11:37:@1176.4]
  assign _T_557 = _T_160 ? 1'h0 : _T_556; // @[Lookup.scala 11:37:@1177.4]
  assign _T_558 = _T_156 ? 1'h0 : _T_557; // @[Lookup.scala 11:37:@1178.4]
  assign _T_559 = _T_152 ? 1'h0 : _T_558; // @[Lookup.scala 11:37:@1179.4]
  assign _T_560 = _T_148 ? 1'h0 : _T_559; // @[Lookup.scala 11:37:@1180.4]
  assign _T_561 = _T_144 ? 1'h0 : _T_560; // @[Lookup.scala 11:37:@1181.4]
  assign _T_562 = _T_140 ? 1'h0 : _T_561; // @[Lookup.scala 11:37:@1182.4]
  assign _T_563 = _T_136 ? 1'h0 : _T_562; // @[Lookup.scala 11:37:@1183.4]
  assign _T_564 = _T_132 ? 1'h0 : _T_563; // @[Lookup.scala 11:37:@1184.4]
  assign _T_565 = _T_128 ? 1'h0 : _T_564; // @[Lookup.scala 11:37:@1185.4]
  assign ctlsig_4 = _T_124 ? 1'h0 : _T_565; // @[Lookup.scala 11:37:@1186.4]
  assign _T_573 = _T_292 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:@1194.4]
  assign _T_574 = _T_288 ? 2'h3 : _T_573; // @[Lookup.scala 11:37:@1195.4]
  assign _T_575 = _T_284 ? 2'h3 : _T_574; // @[Lookup.scala 11:37:@1196.4]
  assign _T_576 = _T_280 ? 2'h3 : _T_575; // @[Lookup.scala 11:37:@1197.4]
  assign _T_577 = _T_276 ? 2'h3 : _T_576; // @[Lookup.scala 11:37:@1198.4]
  assign _T_578 = _T_272 ? 2'h3 : _T_577; // @[Lookup.scala 11:37:@1199.4]
  assign _T_579 = _T_268 ? 2'h0 : _T_578; // @[Lookup.scala 11:37:@1200.4]
  assign _T_580 = _T_264 ? 2'h0 : _T_579; // @[Lookup.scala 11:37:@1201.4]
  assign _T_581 = _T_260 ? 2'h0 : _T_580; // @[Lookup.scala 11:37:@1202.4]
  assign _T_582 = _T_256 ? 2'h0 : _T_581; // @[Lookup.scala 11:37:@1203.4]
  assign _T_583 = _T_252 ? 2'h0 : _T_582; // @[Lookup.scala 11:37:@1204.4]
  assign _T_584 = _T_248 ? 2'h0 : _T_583; // @[Lookup.scala 11:37:@1205.4]
  assign _T_585 = _T_244 ? 2'h0 : _T_584; // @[Lookup.scala 11:37:@1206.4]
  assign _T_586 = _T_240 ? 2'h0 : _T_585; // @[Lookup.scala 11:37:@1207.4]
  assign _T_587 = _T_236 ? 2'h0 : _T_586; // @[Lookup.scala 11:37:@1208.4]
  assign _T_588 = _T_232 ? 2'h0 : _T_587; // @[Lookup.scala 11:37:@1209.4]
  assign _T_589 = _T_228 ? 2'h0 : _T_588; // @[Lookup.scala 11:37:@1210.4]
  assign _T_590 = _T_224 ? 2'h0 : _T_589; // @[Lookup.scala 11:37:@1211.4]
  assign _T_591 = _T_220 ? 2'h0 : _T_590; // @[Lookup.scala 11:37:@1212.4]
  assign _T_592 = _T_216 ? 2'h0 : _T_591; // @[Lookup.scala 11:37:@1213.4]
  assign _T_593 = _T_212 ? 2'h0 : _T_592; // @[Lookup.scala 11:37:@1214.4]
  assign _T_594 = _T_208 ? 2'h0 : _T_593; // @[Lookup.scala 11:37:@1215.4]
  assign _T_595 = _T_204 ? 2'h0 : _T_594; // @[Lookup.scala 11:37:@1216.4]
  assign _T_596 = _T_200 ? 2'h0 : _T_595; // @[Lookup.scala 11:37:@1217.4]
  assign _T_597 = _T_196 ? 2'h0 : _T_596; // @[Lookup.scala 11:37:@1218.4]
  assign _T_598 = _T_192 ? 2'h0 : _T_597; // @[Lookup.scala 11:37:@1219.4]
  assign _T_599 = _T_188 ? 2'h0 : _T_598; // @[Lookup.scala 11:37:@1220.4]
  assign _T_600 = _T_184 ? 2'h0 : _T_599; // @[Lookup.scala 11:37:@1221.4]
  assign _T_601 = _T_180 ? 2'h1 : _T_600; // @[Lookup.scala 11:37:@1222.4]
  assign _T_602 = _T_176 ? 2'h1 : _T_601; // @[Lookup.scala 11:37:@1223.4]
  assign _T_603 = _T_172 ? 2'h1 : _T_602; // @[Lookup.scala 11:37:@1224.4]
  assign _T_604 = _T_168 ? 2'h1 : _T_603; // @[Lookup.scala 11:37:@1225.4]
  assign _T_605 = _T_164 ? 2'h1 : _T_604; // @[Lookup.scala 11:37:@1226.4]
  assign _T_606 = _T_160 ? 2'h0 : _T_605; // @[Lookup.scala 11:37:@1227.4]
  assign _T_607 = _T_156 ? 2'h0 : _T_606; // @[Lookup.scala 11:37:@1228.4]
  assign _T_608 = _T_152 ? 2'h0 : _T_607; // @[Lookup.scala 11:37:@1229.4]
  assign _T_609 = _T_148 ? 2'h0 : _T_608; // @[Lookup.scala 11:37:@1230.4]
  assign _T_610 = _T_144 ? 2'h0 : _T_609; // @[Lookup.scala 11:37:@1231.4]
  assign _T_611 = _T_140 ? 2'h0 : _T_610; // @[Lookup.scala 11:37:@1232.4]
  assign _T_612 = _T_136 ? 2'h2 : _T_611; // @[Lookup.scala 11:37:@1233.4]
  assign _T_613 = _T_132 ? 2'h2 : _T_612; // @[Lookup.scala 11:37:@1234.4]
  assign _T_614 = _T_128 ? 2'h0 : _T_613; // @[Lookup.scala 11:37:@1235.4]
  assign ctlsig_5 = _T_124 ? 2'h0 : _T_614; // @[Lookup.scala 11:37:@1236.4]
  assign _T_648 = _T_188 ? 3'h1 : 3'h2; // @[Lookup.scala 11:37:@1270.4]
  assign _T_649 = _T_184 ? 3'h0 : _T_648; // @[Lookup.scala 11:37:@1271.4]
  assign _T_650 = _T_180 ? 3'h5 : _T_649; // @[Lookup.scala 11:37:@1272.4]
  assign _T_651 = _T_176 ? 3'h4 : _T_650; // @[Lookup.scala 11:37:@1273.4]
  assign _T_652 = _T_172 ? 3'h2 : _T_651; // @[Lookup.scala 11:37:@1274.4]
  assign _T_653 = _T_168 ? 3'h1 : _T_652; // @[Lookup.scala 11:37:@1275.4]
  assign _T_654 = _T_164 ? 3'h0 : _T_653; // @[Lookup.scala 11:37:@1276.4]
  assign _T_655 = _T_160 ? 3'h0 : _T_654; // @[Lookup.scala 11:37:@1277.4]
  assign _T_656 = _T_156 ? 3'h0 : _T_655; // @[Lookup.scala 11:37:@1278.4]
  assign _T_657 = _T_152 ? 3'h0 : _T_656; // @[Lookup.scala 11:37:@1279.4]
  assign _T_658 = _T_148 ? 3'h0 : _T_657; // @[Lookup.scala 11:37:@1280.4]
  assign _T_659 = _T_144 ? 3'h0 : _T_658; // @[Lookup.scala 11:37:@1281.4]
  assign _T_660 = _T_140 ? 3'h0 : _T_659; // @[Lookup.scala 11:37:@1282.4]
  assign _T_661 = _T_136 ? 3'h2 : _T_660; // @[Lookup.scala 11:37:@1283.4]
  assign _T_662 = _T_132 ? 3'h2 : _T_661; // @[Lookup.scala 11:37:@1284.4]
  assign _T_663 = _T_128 ? 3'h2 : _T_662; // @[Lookup.scala 11:37:@1285.4]
  assign ctlsig_6 = _T_124 ? 3'h2 : _T_663; // @[Lookup.scala 11:37:@1286.4]
  assign _T_664 = _T_320 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:@1287.4]
  assign _T_665 = _T_316 ? 2'h0 : _T_664; // @[Lookup.scala 11:37:@1288.4]
  assign _T_666 = _T_312 ? 2'h3 : _T_665; // @[Lookup.scala 11:37:@1289.4]
  assign _T_667 = _T_308 ? 2'h3 : _T_666; // @[Lookup.scala 11:37:@1290.4]
  assign _T_668 = _T_304 ? 2'h3 : _T_667; // @[Lookup.scala 11:37:@1291.4]
  assign _T_669 = _T_300 ? 2'h0 : _T_668; // @[Lookup.scala 11:37:@1292.4]
  assign _T_670 = _T_296 ? 2'h0 : _T_669; // @[Lookup.scala 11:37:@1293.4]
  assign _T_671 = _T_292 ? 2'h0 : _T_670; // @[Lookup.scala 11:37:@1294.4]
  assign _T_672 = _T_288 ? 2'h0 : _T_671; // @[Lookup.scala 11:37:@1295.4]
  assign _T_673 = _T_284 ? 2'h0 : _T_672; // @[Lookup.scala 11:37:@1296.4]
  assign _T_674 = _T_280 ? 2'h0 : _T_673; // @[Lookup.scala 11:37:@1297.4]
  assign _T_675 = _T_276 ? 2'h0 : _T_674; // @[Lookup.scala 11:37:@1298.4]
  assign _T_676 = _T_272 ? 2'h0 : _T_675; // @[Lookup.scala 11:37:@1299.4]
  assign _T_677 = _T_268 ? 2'h0 : _T_676; // @[Lookup.scala 11:37:@1300.4]
  assign _T_678 = _T_264 ? 2'h0 : _T_677; // @[Lookup.scala 11:37:@1301.4]
  assign _T_679 = _T_260 ? 2'h0 : _T_678; // @[Lookup.scala 11:37:@1302.4]
  assign _T_680 = _T_256 ? 2'h0 : _T_679; // @[Lookup.scala 11:37:@1303.4]
  assign _T_681 = _T_252 ? 2'h0 : _T_680; // @[Lookup.scala 11:37:@1304.4]
  assign _T_682 = _T_248 ? 2'h0 : _T_681; // @[Lookup.scala 11:37:@1305.4]
  assign _T_683 = _T_244 ? 2'h0 : _T_682; // @[Lookup.scala 11:37:@1306.4]
  assign _T_684 = _T_240 ? 2'h0 : _T_683; // @[Lookup.scala 11:37:@1307.4]
  assign _T_685 = _T_236 ? 2'h0 : _T_684; // @[Lookup.scala 11:37:@1308.4]
  assign _T_686 = _T_232 ? 2'h0 : _T_685; // @[Lookup.scala 11:37:@1309.4]
  assign _T_687 = _T_228 ? 2'h0 : _T_686; // @[Lookup.scala 11:37:@1310.4]
  assign _T_688 = _T_224 ? 2'h0 : _T_687; // @[Lookup.scala 11:37:@1311.4]
  assign _T_689 = _T_220 ? 2'h0 : _T_688; // @[Lookup.scala 11:37:@1312.4]
  assign _T_690 = _T_216 ? 2'h0 : _T_689; // @[Lookup.scala 11:37:@1313.4]
  assign _T_691 = _T_212 ? 2'h0 : _T_690; // @[Lookup.scala 11:37:@1314.4]
  assign _T_692 = _T_208 ? 2'h0 : _T_691; // @[Lookup.scala 11:37:@1315.4]
  assign _T_693 = _T_204 ? 2'h0 : _T_692; // @[Lookup.scala 11:37:@1316.4]
  assign _T_694 = _T_200 ? 2'h0 : _T_693; // @[Lookup.scala 11:37:@1317.4]
  assign _T_695 = _T_196 ? 2'h0 : _T_694; // @[Lookup.scala 11:37:@1318.4]
  assign _T_696 = _T_192 ? 2'h0 : _T_695; // @[Lookup.scala 11:37:@1319.4]
  assign _T_697 = _T_188 ? 2'h0 : _T_696; // @[Lookup.scala 11:37:@1320.4]
  assign _T_698 = _T_184 ? 2'h0 : _T_697; // @[Lookup.scala 11:37:@1321.4]
  assign _T_699 = _T_180 ? 2'h0 : _T_698; // @[Lookup.scala 11:37:@1322.4]
  assign _T_700 = _T_176 ? 2'h0 : _T_699; // @[Lookup.scala 11:37:@1323.4]
  assign _T_701 = _T_172 ? 2'h0 : _T_700; // @[Lookup.scala 11:37:@1324.4]
  assign _T_702 = _T_168 ? 2'h0 : _T_701; // @[Lookup.scala 11:37:@1325.4]
  assign _T_703 = _T_164 ? 2'h0 : _T_702; // @[Lookup.scala 11:37:@1326.4]
  assign _T_704 = _T_160 ? 2'h1 : _T_703; // @[Lookup.scala 11:37:@1327.4]
  assign _T_705 = _T_156 ? 2'h1 : _T_704; // @[Lookup.scala 11:37:@1328.4]
  assign _T_706 = _T_152 ? 2'h1 : _T_705; // @[Lookup.scala 11:37:@1329.4]
  assign _T_707 = _T_148 ? 2'h1 : _T_706; // @[Lookup.scala 11:37:@1330.4]
  assign _T_708 = _T_144 ? 2'h1 : _T_707; // @[Lookup.scala 11:37:@1331.4]
  assign _T_709 = _T_140 ? 2'h1 : _T_708; // @[Lookup.scala 11:37:@1332.4]
  assign _T_710 = _T_136 ? 2'h2 : _T_709; // @[Lookup.scala 11:37:@1333.4]
  assign _T_711 = _T_132 ? 2'h2 : _T_710; // @[Lookup.scala 11:37:@1334.4]
  assign _T_712 = _T_128 ? 2'h0 : _T_711; // @[Lookup.scala 11:37:@1335.4]
  assign ctlsig_7 = _T_124 ? 2'h0 : _T_712; // @[Lookup.scala 11:37:@1336.4]
  assign _T_753 = _T_160 ? 3'h5 : 3'h7; // @[Lookup.scala 11:37:@1377.4]
  assign _T_754 = _T_156 ? 3'h4 : _T_753; // @[Lookup.scala 11:37:@1378.4]
  assign _T_755 = _T_152 ? 3'h3 : _T_754; // @[Lookup.scala 11:37:@1379.4]
  assign _T_756 = _T_148 ? 3'h2 : _T_755; // @[Lookup.scala 11:37:@1380.4]
  assign _T_757 = _T_144 ? 3'h1 : _T_756; // @[Lookup.scala 11:37:@1381.4]
  assign _T_758 = _T_140 ? 3'h0 : _T_757; // @[Lookup.scala 11:37:@1382.4]
  assign _T_759 = _T_136 ? 3'h7 : _T_758; // @[Lookup.scala 11:37:@1383.4]
  assign _T_760 = _T_132 ? 3'h7 : _T_759; // @[Lookup.scala 11:37:@1384.4]
  assign _T_761 = _T_128 ? 3'h7 : _T_760; // @[Lookup.scala 11:37:@1385.4]
  assign br_sel = _T_124 ? 3'h7 : _T_761; // @[Lookup.scala 11:37:@1386.4]
  assign _T_769 = _T_292 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:@1394.4]
  assign _T_770 = _T_288 ? 2'h2 : _T_769; // @[Lookup.scala 11:37:@1395.4]
  assign _T_771 = _T_284 ? 2'h2 : _T_770; // @[Lookup.scala 11:37:@1396.4]
  assign _T_772 = _T_280 ? 2'h0 : _T_771; // @[Lookup.scala 11:37:@1397.4]
  assign _T_773 = _T_276 ? 2'h0 : _T_772; // @[Lookup.scala 11:37:@1398.4]
  assign _T_774 = _T_272 ? 2'h0 : _T_773; // @[Lookup.scala 11:37:@1399.4]
  assign _T_775 = _T_268 ? 2'h0 : _T_774; // @[Lookup.scala 11:37:@1400.4]
  assign _T_776 = _T_264 ? 2'h0 : _T_775; // @[Lookup.scala 11:37:@1401.4]
  assign _T_777 = _T_260 ? 2'h0 : _T_776; // @[Lookup.scala 11:37:@1402.4]
  assign _T_778 = _T_256 ? 2'h0 : _T_777; // @[Lookup.scala 11:37:@1403.4]
  assign _T_779 = _T_252 ? 2'h0 : _T_778; // @[Lookup.scala 11:37:@1404.4]
  assign _T_780 = _T_248 ? 2'h0 : _T_779; // @[Lookup.scala 11:37:@1405.4]
  assign _T_781 = _T_244 ? 2'h0 : _T_780; // @[Lookup.scala 11:37:@1406.4]
  assign _T_782 = _T_240 ? 2'h0 : _T_781; // @[Lookup.scala 11:37:@1407.4]
  assign _T_783 = _T_236 ? 2'h0 : _T_782; // @[Lookup.scala 11:37:@1408.4]
  assign _T_784 = _T_232 ? 2'h0 : _T_783; // @[Lookup.scala 11:37:@1409.4]
  assign _T_785 = _T_228 ? 2'h0 : _T_784; // @[Lookup.scala 11:37:@1410.4]
  assign _T_786 = _T_224 ? 2'h0 : _T_785; // @[Lookup.scala 11:37:@1411.4]
  assign _T_787 = _T_220 ? 2'h0 : _T_786; // @[Lookup.scala 11:37:@1412.4]
  assign _T_788 = _T_216 ? 2'h0 : _T_787; // @[Lookup.scala 11:37:@1413.4]
  assign _T_789 = _T_212 ? 2'h0 : _T_788; // @[Lookup.scala 11:37:@1414.4]
  assign _T_790 = _T_208 ? 2'h0 : _T_789; // @[Lookup.scala 11:37:@1415.4]
  assign _T_791 = _T_204 ? 2'h0 : _T_790; // @[Lookup.scala 11:37:@1416.4]
  assign _T_792 = _T_200 ? 2'h0 : _T_791; // @[Lookup.scala 11:37:@1417.4]
  assign _T_793 = _T_196 ? 2'h0 : _T_792; // @[Lookup.scala 11:37:@1418.4]
  assign _T_794 = _T_192 ? 2'h0 : _T_793; // @[Lookup.scala 11:37:@1419.4]
  assign _T_795 = _T_188 ? 2'h0 : _T_794; // @[Lookup.scala 11:37:@1420.4]
  assign _T_796 = _T_184 ? 2'h0 : _T_795; // @[Lookup.scala 11:37:@1421.4]
  assign _T_797 = _T_180 ? 2'h0 : _T_796; // @[Lookup.scala 11:37:@1422.4]
  assign _T_798 = _T_176 ? 2'h0 : _T_797; // @[Lookup.scala 11:37:@1423.4]
  assign _T_799 = _T_172 ? 2'h0 : _T_798; // @[Lookup.scala 11:37:@1424.4]
  assign _T_800 = _T_168 ? 2'h0 : _T_799; // @[Lookup.scala 11:37:@1425.4]
  assign _T_801 = _T_164 ? 2'h0 : _T_800; // @[Lookup.scala 11:37:@1426.4]
  assign _T_802 = _T_160 ? 2'h1 : _T_801; // @[Lookup.scala 11:37:@1427.4]
  assign _T_803 = _T_156 ? 2'h1 : _T_802; // @[Lookup.scala 11:37:@1428.4]
  assign _T_804 = _T_152 ? 2'h1 : _T_803; // @[Lookup.scala 11:37:@1429.4]
  assign _T_805 = _T_148 ? 2'h1 : _T_804; // @[Lookup.scala 11:37:@1430.4]
  assign _T_806 = _T_144 ? 2'h1 : _T_805; // @[Lookup.scala 11:37:@1431.4]
  assign _T_807 = _T_140 ? 2'h1 : _T_806; // @[Lookup.scala 11:37:@1432.4]
  assign _T_808 = _T_136 ? 2'h0 : _T_807; // @[Lookup.scala 11:37:@1433.4]
  assign _T_809 = _T_132 ? 2'h1 : _T_808; // @[Lookup.scala 11:37:@1434.4]
  assign _T_810 = _T_128 ? 2'h1 : _T_809; // @[Lookup.scala 11:37:@1435.4]
  assign ctlsig_9 = _T_124 ? 2'h0 : _T_810; // @[Lookup.scala 11:37:@1436.4]
  assign _T_811 = _T_320 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:@1437.4]
  assign _T_812 = _T_316 ? 3'h4 : _T_811; // @[Lookup.scala 11:37:@1438.4]
  assign _T_813 = _T_312 ? 3'h4 : _T_812; // @[Lookup.scala 11:37:@1439.4]
  assign _T_814 = _T_308 ? 3'h4 : _T_813; // @[Lookup.scala 11:37:@1440.4]
  assign _T_815 = _T_304 ? 3'h4 : _T_814; // @[Lookup.scala 11:37:@1441.4]
  assign _T_816 = _T_300 ? 3'h0 : _T_815; // @[Lookup.scala 11:37:@1442.4]
  assign _T_817 = _T_296 ? 3'h0 : _T_816; // @[Lookup.scala 11:37:@1443.4]
  assign _T_818 = _T_292 ? 3'h3 : _T_817; // @[Lookup.scala 11:37:@1444.4]
  assign _T_819 = _T_288 ? 3'h2 : _T_818; // @[Lookup.scala 11:37:@1445.4]
  assign _T_820 = _T_284 ? 3'h1 : _T_819; // @[Lookup.scala 11:37:@1446.4]
  assign _T_821 = _T_280 ? 3'h3 : _T_820; // @[Lookup.scala 11:37:@1447.4]
  assign _T_822 = _T_276 ? 3'h2 : _T_821; // @[Lookup.scala 11:37:@1448.4]
  assign _T_823 = _T_272 ? 3'h1 : _T_822; // @[Lookup.scala 11:37:@1449.4]
  assign _T_824 = _T_268 ? 3'h0 : _T_823; // @[Lookup.scala 11:37:@1450.4]
  assign _T_825 = _T_264 ? 3'h0 : _T_824; // @[Lookup.scala 11:37:@1451.4]
  assign _T_826 = _T_260 ? 3'h0 : _T_825; // @[Lookup.scala 11:37:@1452.4]
  assign _T_827 = _T_256 ? 3'h0 : _T_826; // @[Lookup.scala 11:37:@1453.4]
  assign _T_828 = _T_252 ? 3'h0 : _T_827; // @[Lookup.scala 11:37:@1454.4]
  assign _T_829 = _T_248 ? 3'h0 : _T_828; // @[Lookup.scala 11:37:@1455.4]
  assign _T_830 = _T_244 ? 3'h0 : _T_829; // @[Lookup.scala 11:37:@1456.4]
  assign _T_831 = _T_240 ? 3'h0 : _T_830; // @[Lookup.scala 11:37:@1457.4]
  assign _T_832 = _T_236 ? 3'h0 : _T_831; // @[Lookup.scala 11:37:@1458.4]
  assign _T_833 = _T_232 ? 3'h0 : _T_832; // @[Lookup.scala 11:37:@1459.4]
  assign _T_834 = _T_228 ? 3'h0 : _T_833; // @[Lookup.scala 11:37:@1460.4]
  assign _T_835 = _T_224 ? 3'h0 : _T_834; // @[Lookup.scala 11:37:@1461.4]
  assign _T_836 = _T_220 ? 3'h0 : _T_835; // @[Lookup.scala 11:37:@1462.4]
  assign _T_837 = _T_216 ? 3'h0 : _T_836; // @[Lookup.scala 11:37:@1463.4]
  assign _T_838 = _T_212 ? 3'h0 : _T_837; // @[Lookup.scala 11:37:@1464.4]
  assign _T_839 = _T_208 ? 3'h0 : _T_838; // @[Lookup.scala 11:37:@1465.4]
  assign _T_840 = _T_204 ? 3'h0 : _T_839; // @[Lookup.scala 11:37:@1466.4]
  assign _T_841 = _T_200 ? 3'h0 : _T_840; // @[Lookup.scala 11:37:@1467.4]
  assign _T_842 = _T_196 ? 3'h0 : _T_841; // @[Lookup.scala 11:37:@1468.4]
  assign _T_843 = _T_192 ? 3'h0 : _T_842; // @[Lookup.scala 11:37:@1469.4]
  assign _T_844 = _T_188 ? 3'h0 : _T_843; // @[Lookup.scala 11:37:@1470.4]
  assign _T_845 = _T_184 ? 3'h0 : _T_844; // @[Lookup.scala 11:37:@1471.4]
  assign _T_846 = _T_180 ? 3'h0 : _T_845; // @[Lookup.scala 11:37:@1472.4]
  assign _T_847 = _T_176 ? 3'h0 : _T_846; // @[Lookup.scala 11:37:@1473.4]
  assign _T_848 = _T_172 ? 3'h0 : _T_847; // @[Lookup.scala 11:37:@1474.4]
  assign _T_849 = _T_168 ? 3'h0 : _T_848; // @[Lookup.scala 11:37:@1475.4]
  assign _T_850 = _T_164 ? 3'h0 : _T_849; // @[Lookup.scala 11:37:@1476.4]
  assign _T_851 = _T_160 ? 3'h0 : _T_850; // @[Lookup.scala 11:37:@1477.4]
  assign _T_852 = _T_156 ? 3'h0 : _T_851; // @[Lookup.scala 11:37:@1478.4]
  assign _T_853 = _T_152 ? 3'h0 : _T_852; // @[Lookup.scala 11:37:@1479.4]
  assign _T_854 = _T_148 ? 3'h0 : _T_853; // @[Lookup.scala 11:37:@1480.4]
  assign _T_855 = _T_144 ? 3'h0 : _T_854; // @[Lookup.scala 11:37:@1481.4]
  assign _T_856 = _T_140 ? 3'h0 : _T_855; // @[Lookup.scala 11:37:@1482.4]
  assign _T_857 = _T_136 ? 3'h0 : _T_856; // @[Lookup.scala 11:37:@1483.4]
  assign _T_858 = _T_132 ? 3'h0 : _T_857; // @[Lookup.scala 11:37:@1484.4]
  assign _T_859 = _T_128 ? 3'h0 : _T_858; // @[Lookup.scala 11:37:@1485.4]
  assign csr_cmd = _T_124 ? 3'h0 : _T_859; // @[Lookup.scala 11:37:@1486.4]
  assign _T_861 = _T_316 ? 1'h1 : _T_320; // @[Lookup.scala 11:37:@1488.4]
  assign _T_862 = _T_312 ? 1'h1 : _T_861; // @[Lookup.scala 11:37:@1489.4]
  assign _T_863 = _T_308 ? 1'h1 : _T_862; // @[Lookup.scala 11:37:@1490.4]
  assign _T_864 = _T_304 ? 1'h1 : _T_863; // @[Lookup.scala 11:37:@1491.4]
  assign _T_865 = _T_300 ? 1'h1 : _T_864; // @[Lookup.scala 11:37:@1492.4]
  assign _T_866 = _T_296 ? 1'h1 : _T_865; // @[Lookup.scala 11:37:@1493.4]
  assign _T_867 = _T_292 ? 1'h1 : _T_866; // @[Lookup.scala 11:37:@1494.4]
  assign _T_868 = _T_288 ? 1'h1 : _T_867; // @[Lookup.scala 11:37:@1495.4]
  assign _T_869 = _T_284 ? 1'h1 : _T_868; // @[Lookup.scala 11:37:@1496.4]
  assign _T_870 = _T_280 ? 1'h1 : _T_869; // @[Lookup.scala 11:37:@1497.4]
  assign _T_871 = _T_276 ? 1'h1 : _T_870; // @[Lookup.scala 11:37:@1498.4]
  assign _T_872 = _T_272 ? 1'h1 : _T_871; // @[Lookup.scala 11:37:@1499.4]
  assign _T_873 = _T_268 ? 1'h1 : _T_872; // @[Lookup.scala 11:37:@1500.4]
  assign _T_874 = _T_264 ? 1'h1 : _T_873; // @[Lookup.scala 11:37:@1501.4]
  assign _T_875 = _T_260 ? 1'h1 : _T_874; // @[Lookup.scala 11:37:@1502.4]
  assign _T_876 = _T_256 ? 1'h1 : _T_875; // @[Lookup.scala 11:37:@1503.4]
  assign _T_877 = _T_252 ? 1'h1 : _T_876; // @[Lookup.scala 11:37:@1504.4]
  assign _T_878 = _T_248 ? 1'h1 : _T_877; // @[Lookup.scala 11:37:@1505.4]
  assign _T_879 = _T_244 ? 1'h1 : _T_878; // @[Lookup.scala 11:37:@1506.4]
  assign _T_880 = _T_240 ? 1'h1 : _T_879; // @[Lookup.scala 11:37:@1507.4]
  assign _T_881 = _T_236 ? 1'h1 : _T_880; // @[Lookup.scala 11:37:@1508.4]
  assign _T_882 = _T_232 ? 1'h1 : _T_881; // @[Lookup.scala 11:37:@1509.4]
  assign _T_883 = _T_228 ? 1'h1 : _T_882; // @[Lookup.scala 11:37:@1510.4]
  assign _T_884 = _T_224 ? 1'h1 : _T_883; // @[Lookup.scala 11:37:@1511.4]
  assign _T_885 = _T_220 ? 1'h1 : _T_884; // @[Lookup.scala 11:37:@1512.4]
  assign _T_886 = _T_216 ? 1'h1 : _T_885; // @[Lookup.scala 11:37:@1513.4]
  assign _T_887 = _T_212 ? 1'h1 : _T_886; // @[Lookup.scala 11:37:@1514.4]
  assign _T_888 = _T_208 ? 1'h1 : _T_887; // @[Lookup.scala 11:37:@1515.4]
  assign _T_889 = _T_204 ? 1'h1 : _T_888; // @[Lookup.scala 11:37:@1516.4]
  assign _T_890 = _T_200 ? 1'h1 : _T_889; // @[Lookup.scala 11:37:@1517.4]
  assign _T_891 = _T_196 ? 1'h1 : _T_890; // @[Lookup.scala 11:37:@1518.4]
  assign _T_892 = _T_192 ? 1'h1 : _T_891; // @[Lookup.scala 11:37:@1519.4]
  assign _T_893 = _T_188 ? 1'h1 : _T_892; // @[Lookup.scala 11:37:@1520.4]
  assign _T_894 = _T_184 ? 1'h1 : _T_893; // @[Lookup.scala 11:37:@1521.4]
  assign _T_895 = _T_180 ? 1'h1 : _T_894; // @[Lookup.scala 11:37:@1522.4]
  assign _T_896 = _T_176 ? 1'h1 : _T_895; // @[Lookup.scala 11:37:@1523.4]
  assign _T_897 = _T_172 ? 1'h1 : _T_896; // @[Lookup.scala 11:37:@1524.4]
  assign _T_898 = _T_168 ? 1'h1 : _T_897; // @[Lookup.scala 11:37:@1525.4]
  assign _T_899 = _T_164 ? 1'h1 : _T_898; // @[Lookup.scala 11:37:@1526.4]
  assign _T_900 = _T_160 ? 1'h1 : _T_899; // @[Lookup.scala 11:37:@1527.4]
  assign _T_901 = _T_156 ? 1'h1 : _T_900; // @[Lookup.scala 11:37:@1528.4]
  assign _T_902 = _T_152 ? 1'h1 : _T_901; // @[Lookup.scala 11:37:@1529.4]
  assign _T_903 = _T_148 ? 1'h1 : _T_902; // @[Lookup.scala 11:37:@1530.4]
  assign _T_904 = _T_144 ? 1'h1 : _T_903; // @[Lookup.scala 11:37:@1531.4]
  assign _T_905 = _T_140 ? 1'h1 : _T_904; // @[Lookup.scala 11:37:@1532.4]
  assign _T_906 = _T_136 ? 1'h1 : _T_905; // @[Lookup.scala 11:37:@1533.4]
  assign _T_907 = _T_132 ? 1'h1 : _T_906; // @[Lookup.scala 11:37:@1534.4]
  assign _T_908 = _T_128 ? 1'h1 : _T_907; // @[Lookup.scala 11:37:@1535.4]
  assign ctlsig_11 = _T_124 ? 1'h1 : _T_908; // @[Lookup.scala 11:37:@1536.4]
  assign _T_909 = io_c2d_cexcp | io_d2c_dexcp; // @[rvcpath.scala 134:39:@1544.4]
  assign _T_910 = _T_909 ? 2'h3 : ctlsig_7; // @[rvcpath.scala 134:25:@1545.4]
  assign _T_911 = ctlsig_11 == 1'h0; // @[rvcpath.scala 139:33:@1550.4]
  assign _T_913 = io_c2d_cexcp ? 4'h2 : 4'h0; // @[rvcpath.scala 140:25:@1552.4]
  assign io_c2d_alu_func = alu_func;
  assign io_c2d_op2_sel = ctlsig_1;
  assign io_c2d_reg_wren = ctlsig_2;
  assign io_c2d_mem_wren = ctlsig_3;
  assign io_c2d_mem_en = ctlsig_4;
  assign io_c2d_wb_sel = ctlsig_5;
  assign io_c2d_mem_type = ctlsig_6;
  assign io_c2d_pc_sel = _T_910;
  assign io_c2d_br_sel = br_sel;
  assign io_c2d_op1_sel = ctlsig_9;
  assign io_c2d_csr_cmd = csr_cmd;
  assign io_c2d_cexcp = _T_911;
  assign io_c2d_ccause = _T_913;
endmodule
module rvcsr( // @[:@1555.2]
  input         clock, // @[:@1556.4]
  input         reset, // @[:@1557.4]
  input  [11:0] io_addr, // @[:@1558.4]
  input  [31:0] io_wdata, // @[:@1558.4]
  output [31:0] io_rdata, // @[:@1558.4]
  input  [2:0]  io_op, // @[:@1558.4]
  input  [31:0] io_core_pc, // @[:@1558.4]
  input         io_core_excp, // @[:@1558.4]
  input  [3:0]  io_core_cause, // @[:@1558.4]
  output        io_csr_excp, // @[:@1558.4]
  output [31:0] io_csr_evec // @[:@1558.4]
);
  reg [1:0] reg_priv; // @[rvcsr.scala 186:23:@1570.4]
  reg [31:0] _RAND_0;
  reg [31:0] reg_mstatus; // @[rvcsr.scala 188:26:@1571.4]
  reg [31:0] _RAND_1;
  reg [31:0] reg_mtvec; // @[rvcsr.scala 189:24:@1572.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_medeleg; // @[rvcsr.scala 190:26:@1573.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_mideleg; // @[rvcsr.scala 191:26:@1574.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_mip; // @[rvcsr.scala 192:22:@1575.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_mie; // @[rvcsr.scala 193:22:@1576.4]
  reg [31:0] _RAND_6;
  reg [63:0] reg_mtime; // @[rvcsr.scala 194:24:@1577.4]
  reg [63:0] _RAND_7;
  reg [63:0] reg_mtimecmp; // @[rvcsr.scala 196:27:@1578.4]
  reg [63:0] _RAND_8;
  reg [63:0] reg_mcycle; // @[rvcsr.scala 197:25:@1579.4]
  reg [63:0] _RAND_9;
  reg [63:0] reg_minstret; // @[rvcsr.scala 198:27:@1580.4]
  reg [63:0] _RAND_10;
  reg [63:0] reg_mhpmcounters_0; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_11;
  reg [63:0] reg_mhpmcounters_1; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_12;
  reg [63:0] reg_mhpmcounters_2; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_13;
  reg [63:0] reg_mhpmcounters_3; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_14;
  reg [63:0] reg_mhpmcounters_4; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_15;
  reg [63:0] reg_mhpmcounters_5; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_16;
  reg [63:0] reg_mhpmcounters_6; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_17;
  reg [63:0] reg_mhpmcounters_7; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_18;
  reg [63:0] reg_mhpmcounters_8; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_19;
  reg [63:0] reg_mhpmcounters_9; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_20;
  reg [63:0] reg_mhpmcounters_10; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_21;
  reg [63:0] reg_mhpmcounters_11; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_22;
  reg [63:0] reg_mhpmcounters_12; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_23;
  reg [63:0] reg_mhpmcounters_13; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_24;
  reg [63:0] reg_mhpmcounters_14; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_25;
  reg [63:0] reg_mhpmcounters_15; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_26;
  reg [63:0] reg_mhpmcounters_16; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_27;
  reg [63:0] reg_mhpmcounters_17; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_28;
  reg [63:0] reg_mhpmcounters_18; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_29;
  reg [63:0] reg_mhpmcounters_19; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_30;
  reg [63:0] reg_mhpmcounters_20; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_31;
  reg [63:0] reg_mhpmcounters_21; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_32;
  reg [63:0] reg_mhpmcounters_22; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_33;
  reg [63:0] reg_mhpmcounters_23; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_34;
  reg [63:0] reg_mhpmcounters_24; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_35;
  reg [63:0] reg_mhpmcounters_25; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_36;
  reg [63:0] reg_mhpmcounters_26; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_37;
  reg [63:0] reg_mhpmcounters_27; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_38;
  reg [63:0] reg_mhpmcounters_28; // @[rvcsr.scala 200:31:@1581.4]
  reg [63:0] _RAND_39;
  reg [31:0] reg_mhpmevents_0; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_40;
  reg [31:0] reg_mhpmevents_1; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_41;
  reg [31:0] reg_mhpmevents_2; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_42;
  reg [31:0] reg_mhpmevents_3; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_43;
  reg [31:0] reg_mhpmevents_4; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_44;
  reg [31:0] reg_mhpmevents_5; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_45;
  reg [31:0] reg_mhpmevents_6; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_46;
  reg [31:0] reg_mhpmevents_7; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_47;
  reg [31:0] reg_mhpmevents_8; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_48;
  reg [31:0] reg_mhpmevents_9; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_49;
  reg [31:0] reg_mhpmevents_10; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_50;
  reg [31:0] reg_mhpmevents_11; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_51;
  reg [31:0] reg_mhpmevents_12; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_52;
  reg [31:0] reg_mhpmevents_13; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_53;
  reg [31:0] reg_mhpmevents_14; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_54;
  reg [31:0] reg_mhpmevents_15; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_55;
  reg [31:0] reg_mhpmevents_16; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_56;
  reg [31:0] reg_mhpmevents_17; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_57;
  reg [31:0] reg_mhpmevents_18; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_58;
  reg [31:0] reg_mhpmevents_19; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_59;
  reg [31:0] reg_mhpmevents_20; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_60;
  reg [31:0] reg_mhpmevents_21; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_61;
  reg [31:0] reg_mhpmevents_22; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_62;
  reg [31:0] reg_mhpmevents_23; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_63;
  reg [31:0] reg_mhpmevents_24; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_64;
  reg [31:0] reg_mhpmevents_25; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_65;
  reg [31:0] reg_mhpmevents_26; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_66;
  reg [31:0] reg_mhpmevents_27; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_67;
  reg [31:0] reg_mhpmevents_28; // @[rvcsr.scala 201:29:@1582.4]
  reg [31:0] _RAND_68;
  reg [31:0] reg_mcounteren; // @[rvcsr.scala 203:29:@1583.4]
  reg [31:0] _RAND_69;
  reg [31:0] reg_mscratch; // @[rvcsr.scala 204:27:@1584.4]
  reg [31:0] _RAND_70;
  reg [31:0] reg_mepc; // @[rvcsr.scala 205:23:@1585.4]
  reg [31:0] _RAND_71;
  reg [31:0] reg_mcause; // @[rvcsr.scala 206:25:@1586.4]
  reg [31:0] _RAND_72;
  reg [31:0] reg_mtval; // @[rvcsr.scala 207:24:@1587.4]
  reg [31:0] _RAND_73;
  reg [31:0] reg_dcsr; // @[rvcsr.scala 211:23:@1589.4]
  reg [31:0] _RAND_74;
  reg [31:0] reg_dpc; // @[rvcsr.scala 212:22:@1590.4]
  reg [31:0] _RAND_75;
  reg [31:0] reg_dscratch0; // @[rvcsr.scala 213:28:@1591.4]
  reg [31:0] _RAND_76;
  reg [31:0] reg_dscratch1; // @[rvcsr.scala 214:28:@1592.4]
  reg [31:0] _RAND_77;
  wire [31:0] _T_107; // @[rvcsr.scala 253:38:@1594.4]
  wire [31:0] _T_108; // @[rvcsr.scala 254:42:@1595.4]
  wire [31:0] _T_111; // @[rvcsr.scala 258:36:@1598.4]
  wire [31:0] _T_112; // @[rvcsr.scala 259:42:@1599.4]
  wire [31:0] _T_113; // @[rvcsr.scala 260:37:@1600.4]
  wire [31:0] _T_115; // @[rvcsr.scala 273:73:@1602.4]
  wire [31:0] _T_116; // @[rvcsr.scala 274:74:@1603.4]
  wire [31:0] _T_117; // @[rvcsr.scala 273:73:@1604.4]
  wire [31:0] _T_118; // @[rvcsr.scala 274:74:@1605.4]
  wire [31:0] _T_119; // @[rvcsr.scala 273:73:@1606.4]
  wire [31:0] _T_120; // @[rvcsr.scala 274:74:@1607.4]
  wire [31:0] _T_121; // @[rvcsr.scala 273:73:@1608.4]
  wire [31:0] _T_122; // @[rvcsr.scala 274:74:@1609.4]
  wire [31:0] _T_123; // @[rvcsr.scala 273:73:@1610.4]
  wire [31:0] _T_124; // @[rvcsr.scala 274:74:@1611.4]
  wire [31:0] _T_125; // @[rvcsr.scala 273:73:@1612.4]
  wire [31:0] _T_126; // @[rvcsr.scala 274:74:@1613.4]
  wire [31:0] _T_127; // @[rvcsr.scala 273:73:@1614.4]
  wire [31:0] _T_128; // @[rvcsr.scala 274:74:@1615.4]
  wire [31:0] _T_129; // @[rvcsr.scala 273:73:@1616.4]
  wire [31:0] _T_130; // @[rvcsr.scala 274:74:@1617.4]
  wire [31:0] _T_131; // @[rvcsr.scala 273:73:@1618.4]
  wire [31:0] _T_132; // @[rvcsr.scala 274:74:@1619.4]
  wire [31:0] _T_133; // @[rvcsr.scala 273:73:@1620.4]
  wire [31:0] _T_134; // @[rvcsr.scala 274:74:@1621.4]
  wire [31:0] _T_135; // @[rvcsr.scala 273:73:@1622.4]
  wire [31:0] _T_136; // @[rvcsr.scala 274:74:@1623.4]
  wire [31:0] _T_137; // @[rvcsr.scala 273:73:@1624.4]
  wire [31:0] _T_138; // @[rvcsr.scala 274:74:@1625.4]
  wire [31:0] _T_139; // @[rvcsr.scala 273:73:@1626.4]
  wire [31:0] _T_140; // @[rvcsr.scala 274:74:@1627.4]
  wire [31:0] _T_141; // @[rvcsr.scala 273:73:@1628.4]
  wire [31:0] _T_142; // @[rvcsr.scala 274:74:@1629.4]
  wire [31:0] _T_143; // @[rvcsr.scala 273:73:@1630.4]
  wire [31:0] _T_144; // @[rvcsr.scala 274:74:@1631.4]
  wire [31:0] _T_145; // @[rvcsr.scala 273:73:@1632.4]
  wire [31:0] _T_146; // @[rvcsr.scala 274:74:@1633.4]
  wire [31:0] _T_147; // @[rvcsr.scala 273:73:@1634.4]
  wire [31:0] _T_148; // @[rvcsr.scala 274:74:@1635.4]
  wire [31:0] _T_149; // @[rvcsr.scala 273:73:@1636.4]
  wire [31:0] _T_150; // @[rvcsr.scala 274:74:@1637.4]
  wire [31:0] _T_151; // @[rvcsr.scala 273:73:@1638.4]
  wire [31:0] _T_152; // @[rvcsr.scala 274:74:@1639.4]
  wire [31:0] _T_153; // @[rvcsr.scala 273:73:@1640.4]
  wire [31:0] _T_154; // @[rvcsr.scala 274:74:@1641.4]
  wire [31:0] _T_155; // @[rvcsr.scala 273:73:@1642.4]
  wire [31:0] _T_156; // @[rvcsr.scala 274:74:@1643.4]
  wire [31:0] _T_157; // @[rvcsr.scala 273:73:@1644.4]
  wire [31:0] _T_158; // @[rvcsr.scala 274:74:@1645.4]
  wire [31:0] _T_159; // @[rvcsr.scala 273:73:@1646.4]
  wire [31:0] _T_160; // @[rvcsr.scala 274:74:@1647.4]
  wire [31:0] _T_161; // @[rvcsr.scala 273:73:@1648.4]
  wire [31:0] _T_162; // @[rvcsr.scala 274:74:@1649.4]
  wire [31:0] _T_163; // @[rvcsr.scala 273:73:@1650.4]
  wire [31:0] _T_164; // @[rvcsr.scala 274:74:@1651.4]
  wire [31:0] _T_165; // @[rvcsr.scala 273:73:@1652.4]
  wire [31:0] _T_166; // @[rvcsr.scala 274:74:@1653.4]
  wire [31:0] _T_167; // @[rvcsr.scala 273:73:@1654.4]
  wire [31:0] _T_168; // @[rvcsr.scala 274:74:@1655.4]
  wire [31:0] _T_169; // @[rvcsr.scala 273:73:@1656.4]
  wire [31:0] _T_170; // @[rvcsr.scala 274:74:@1657.4]
  wire [31:0] _T_171; // @[rvcsr.scala 273:73:@1658.4]
  wire [31:0] _T_172; // @[rvcsr.scala 274:74:@1659.4]
  wire  counteren_CY; // @[rvcsr.scala 281:48:@1663.4]
  wire  counteren_TM; // @[rvcsr.scala 281:48:@1665.4]
  wire  counteren_IR; // @[rvcsr.scala 281:48:@1667.4]
  wire  counteren_HPM_0; // @[rvcsr.scala 281:48:@1669.4]
  wire  counteren_HPM_1; // @[rvcsr.scala 281:48:@1671.4]
  wire  counteren_HPM_2; // @[rvcsr.scala 281:48:@1673.4]
  wire  counteren_HPM_3; // @[rvcsr.scala 281:48:@1675.4]
  wire  counteren_HPM_4; // @[rvcsr.scala 281:48:@1677.4]
  wire  counteren_HPM_5; // @[rvcsr.scala 281:48:@1679.4]
  wire  counteren_HPM_6; // @[rvcsr.scala 281:48:@1681.4]
  wire  counteren_HPM_7; // @[rvcsr.scala 281:48:@1683.4]
  wire  counteren_HPM_8; // @[rvcsr.scala 281:48:@1685.4]
  wire  counteren_HPM_9; // @[rvcsr.scala 281:48:@1687.4]
  wire  counteren_HPM_10; // @[rvcsr.scala 281:48:@1689.4]
  wire  counteren_HPM_11; // @[rvcsr.scala 281:48:@1691.4]
  wire  counteren_HPM_12; // @[rvcsr.scala 281:48:@1693.4]
  wire  counteren_HPM_13; // @[rvcsr.scala 281:48:@1695.4]
  wire  counteren_HPM_14; // @[rvcsr.scala 281:48:@1697.4]
  wire  counteren_HPM_15; // @[rvcsr.scala 281:48:@1699.4]
  wire  counteren_HPM_16; // @[rvcsr.scala 281:48:@1701.4]
  wire  counteren_HPM_17; // @[rvcsr.scala 281:48:@1703.4]
  wire  counteren_HPM_18; // @[rvcsr.scala 281:48:@1705.4]
  wire  counteren_HPM_19; // @[rvcsr.scala 281:48:@1707.4]
  wire  counteren_HPM_20; // @[rvcsr.scala 281:48:@1709.4]
  wire  counteren_HPM_21; // @[rvcsr.scala 281:48:@1711.4]
  wire  counteren_HPM_22; // @[rvcsr.scala 281:48:@1713.4]
  wire  counteren_HPM_23; // @[rvcsr.scala 281:48:@1715.4]
  wire  counteren_HPM_24; // @[rvcsr.scala 281:48:@1717.4]
  wire  counteren_HPM_25; // @[rvcsr.scala 281:48:@1719.4]
  wire  counteren_HPM_26; // @[rvcsr.scala 281:48:@1721.4]
  wire  counteren_HPM_27; // @[rvcsr.scala 281:48:@1723.4]
  wire  counteren_HPM_28; // @[rvcsr.scala 281:48:@1725.4]
  wire [64:0] _T_216; // @[rvcsr.scala 284:34:@1728.6]
  wire [63:0] _T_217; // @[rvcsr.scala 284:34:@1729.6]
  wire [63:0] _GEN_0; // @[rvcsr.scala 283:24:@1727.4]
  wire [64:0] _T_219; // @[rvcsr.scala 288:32:@1733.6]
  wire [63:0] _T_220; // @[rvcsr.scala 288:32:@1734.6]
  wire [63:0] _GEN_1; // @[rvcsr.scala 287:24:@1732.4]
  wire [64:0] _T_222; // @[rvcsr.scala 292:38:@1738.6]
  wire [63:0] _T_223; // @[rvcsr.scala 292:38:@1739.6]
  wire [63:0] _GEN_2; // @[rvcsr.scala 291:24:@1737.4]
  wire [64:0] _T_225; // @[rvcsr.scala 297:56:@1743.6]
  wire [63:0] _T_226; // @[rvcsr.scala 297:56:@1744.6]
  wire [63:0] _GEN_3; // @[rvcsr.scala 296:32:@1742.4]
  wire [64:0] _T_228; // @[rvcsr.scala 297:56:@1748.6]
  wire [63:0] _T_229; // @[rvcsr.scala 297:56:@1749.6]
  wire [63:0] _GEN_4; // @[rvcsr.scala 296:32:@1747.4]
  wire [64:0] _T_231; // @[rvcsr.scala 297:56:@1753.6]
  wire [63:0] _T_232; // @[rvcsr.scala 297:56:@1754.6]
  wire [63:0] _GEN_5; // @[rvcsr.scala 296:32:@1752.4]
  wire [64:0] _T_234; // @[rvcsr.scala 297:56:@1758.6]
  wire [63:0] _T_235; // @[rvcsr.scala 297:56:@1759.6]
  wire [63:0] _GEN_6; // @[rvcsr.scala 296:32:@1757.4]
  wire [64:0] _T_237; // @[rvcsr.scala 297:56:@1763.6]
  wire [63:0] _T_238; // @[rvcsr.scala 297:56:@1764.6]
  wire [63:0] _GEN_7; // @[rvcsr.scala 296:32:@1762.4]
  wire [64:0] _T_240; // @[rvcsr.scala 297:56:@1768.6]
  wire [63:0] _T_241; // @[rvcsr.scala 297:56:@1769.6]
  wire [63:0] _GEN_8; // @[rvcsr.scala 296:32:@1767.4]
  wire [64:0] _T_243; // @[rvcsr.scala 297:56:@1773.6]
  wire [63:0] _T_244; // @[rvcsr.scala 297:56:@1774.6]
  wire [63:0] _GEN_9; // @[rvcsr.scala 296:32:@1772.4]
  wire [64:0] _T_246; // @[rvcsr.scala 297:56:@1778.6]
  wire [63:0] _T_247; // @[rvcsr.scala 297:56:@1779.6]
  wire [63:0] _GEN_10; // @[rvcsr.scala 296:32:@1777.4]
  wire [64:0] _T_249; // @[rvcsr.scala 297:56:@1783.6]
  wire [63:0] _T_250; // @[rvcsr.scala 297:56:@1784.6]
  wire [63:0] _GEN_11; // @[rvcsr.scala 296:32:@1782.4]
  wire [64:0] _T_252; // @[rvcsr.scala 297:56:@1788.6]
  wire [63:0] _T_253; // @[rvcsr.scala 297:56:@1789.6]
  wire [63:0] _GEN_12; // @[rvcsr.scala 296:32:@1787.4]
  wire [64:0] _T_255; // @[rvcsr.scala 297:56:@1793.6]
  wire [63:0] _T_256; // @[rvcsr.scala 297:56:@1794.6]
  wire [63:0] _GEN_13; // @[rvcsr.scala 296:32:@1792.4]
  wire [64:0] _T_258; // @[rvcsr.scala 297:56:@1798.6]
  wire [63:0] _T_259; // @[rvcsr.scala 297:56:@1799.6]
  wire [63:0] _GEN_14; // @[rvcsr.scala 296:32:@1797.4]
  wire [64:0] _T_261; // @[rvcsr.scala 297:56:@1803.6]
  wire [63:0] _T_262; // @[rvcsr.scala 297:56:@1804.6]
  wire [63:0] _GEN_15; // @[rvcsr.scala 296:32:@1802.4]
  wire [64:0] _T_264; // @[rvcsr.scala 297:56:@1808.6]
  wire [63:0] _T_265; // @[rvcsr.scala 297:56:@1809.6]
  wire [63:0] _GEN_16; // @[rvcsr.scala 296:32:@1807.4]
  wire [64:0] _T_267; // @[rvcsr.scala 297:56:@1813.6]
  wire [63:0] _T_268; // @[rvcsr.scala 297:56:@1814.6]
  wire [63:0] _GEN_17; // @[rvcsr.scala 296:32:@1812.4]
  wire [64:0] _T_270; // @[rvcsr.scala 297:56:@1818.6]
  wire [63:0] _T_271; // @[rvcsr.scala 297:56:@1819.6]
  wire [63:0] _GEN_18; // @[rvcsr.scala 296:32:@1817.4]
  wire [64:0] _T_273; // @[rvcsr.scala 297:56:@1823.6]
  wire [63:0] _T_274; // @[rvcsr.scala 297:56:@1824.6]
  wire [63:0] _GEN_19; // @[rvcsr.scala 296:32:@1822.4]
  wire [64:0] _T_276; // @[rvcsr.scala 297:56:@1828.6]
  wire [63:0] _T_277; // @[rvcsr.scala 297:56:@1829.6]
  wire [63:0] _GEN_20; // @[rvcsr.scala 296:32:@1827.4]
  wire [64:0] _T_279; // @[rvcsr.scala 297:56:@1833.6]
  wire [63:0] _T_280; // @[rvcsr.scala 297:56:@1834.6]
  wire [63:0] _GEN_21; // @[rvcsr.scala 296:32:@1832.4]
  wire [64:0] _T_282; // @[rvcsr.scala 297:56:@1838.6]
  wire [63:0] _T_283; // @[rvcsr.scala 297:56:@1839.6]
  wire [63:0] _GEN_22; // @[rvcsr.scala 296:32:@1837.4]
  wire [64:0] _T_285; // @[rvcsr.scala 297:56:@1843.6]
  wire [63:0] _T_286; // @[rvcsr.scala 297:56:@1844.6]
  wire [63:0] _GEN_23; // @[rvcsr.scala 296:32:@1842.4]
  wire [64:0] _T_288; // @[rvcsr.scala 297:56:@1848.6]
  wire [63:0] _T_289; // @[rvcsr.scala 297:56:@1849.6]
  wire [63:0] _GEN_24; // @[rvcsr.scala 296:32:@1847.4]
  wire [64:0] _T_291; // @[rvcsr.scala 297:56:@1853.6]
  wire [63:0] _T_292; // @[rvcsr.scala 297:56:@1854.6]
  wire [63:0] _GEN_25; // @[rvcsr.scala 296:32:@1852.4]
  wire [64:0] _T_294; // @[rvcsr.scala 297:56:@1858.6]
  wire [63:0] _T_295; // @[rvcsr.scala 297:56:@1859.6]
  wire [63:0] _GEN_26; // @[rvcsr.scala 296:32:@1857.4]
  wire [64:0] _T_297; // @[rvcsr.scala 297:56:@1863.6]
  wire [63:0] _T_298; // @[rvcsr.scala 297:56:@1864.6]
  wire [63:0] _GEN_27; // @[rvcsr.scala 296:32:@1862.4]
  wire [64:0] _T_300; // @[rvcsr.scala 297:56:@1868.6]
  wire [63:0] _T_301; // @[rvcsr.scala 297:56:@1869.6]
  wire [63:0] _GEN_28; // @[rvcsr.scala 296:32:@1867.4]
  wire [64:0] _T_303; // @[rvcsr.scala 297:56:@1873.6]
  wire [63:0] _T_304; // @[rvcsr.scala 297:56:@1874.6]
  wire [63:0] _GEN_29; // @[rvcsr.scala 296:32:@1872.4]
  wire [64:0] _T_306; // @[rvcsr.scala 297:56:@1878.6]
  wire [63:0] _T_307; // @[rvcsr.scala 297:56:@1879.6]
  wire [63:0] _GEN_30; // @[rvcsr.scala 296:32:@1877.4]
  wire [64:0] _T_309; // @[rvcsr.scala 297:56:@1883.6]
  wire [63:0] _T_310; // @[rvcsr.scala 297:56:@1884.6]
  wire [63:0] _GEN_31; // @[rvcsr.scala 296:32:@1882.4]
  wire  _T_318; // @[rvcsr.scala 311:40:@1893.4]
  wire  _T_319; // @[rvcsr.scala 311:40:@1895.4]
  wire  _T_320; // @[rvcsr.scala 311:40:@1897.4]
  wire  _T_321; // @[rvcsr.scala 311:40:@1899.4]
  wire  _T_322; // @[rvcsr.scala 311:40:@1901.4]
  wire  _T_323; // @[rvcsr.scala 311:40:@1903.4]
  wire  _T_324; // @[rvcsr.scala 311:40:@1905.4]
  wire  _T_325; // @[rvcsr.scala 311:40:@1907.4]
  wire  _T_326; // @[rvcsr.scala 311:40:@1909.4]
  wire [1:0] _T_327; // @[rvcsr.scala 311:40:@1911.4]
  wire [1:0] _T_328; // @[rvcsr.scala 311:40:@1913.4]
  wire [1:0] _T_329; // @[rvcsr.scala 311:40:@1915.4]
  wire [1:0] _T_330; // @[rvcsr.scala 311:40:@1917.4]
  wire  _T_331; // @[rvcsr.scala 311:40:@1919.4]
  wire  _T_332; // @[rvcsr.scala 311:40:@1921.4]
  wire  _T_333; // @[rvcsr.scala 311:40:@1923.4]
  wire  _T_334; // @[rvcsr.scala 311:40:@1925.4]
  wire  _T_335; // @[rvcsr.scala 311:40:@1927.4]
  wire  _T_336; // @[rvcsr.scala 311:40:@1929.4]
  wire [7:0] _T_337; // @[rvcsr.scala 311:40:@1931.4]
  wire  _T_338; // @[rvcsr.scala 311:40:@1933.4]
  wire [30:0] _T_344; // @[:@1958.4]
  wire  mie_USIE; // @[rvcsr.scala 313:32:@1960.4]
  wire  mie_SSIE; // @[rvcsr.scala 313:32:@1962.4]
  wire  mie_rsrvd4; // @[rvcsr.scala 313:32:@1964.4]
  wire  _T_348; // @[rvcsr.scala 313:32:@1966.4]
  wire  mie_UTIE; // @[rvcsr.scala 313:32:@1968.4]
  wire  mie_STIE; // @[rvcsr.scala 313:32:@1970.4]
  wire  mie_rsrvd3; // @[rvcsr.scala 313:32:@1972.4]
  wire  _T_352; // @[rvcsr.scala 313:32:@1974.4]
  wire  mie_UEIE; // @[rvcsr.scala 313:32:@1976.4]
  wire  mie_SEIE; // @[rvcsr.scala 313:32:@1978.4]
  wire  mie_rsrvd2; // @[rvcsr.scala 313:32:@1980.4]
  wire  mie_MEIE; // @[rvcsr.scala 313:32:@1982.4]
  wire [18:0] mie_rsrvd1; // @[rvcsr.scala 313:32:@1984.4]
  wire [30:0] _T_363; // @[:@2001.4]
  wire  mip_USIP; // @[rvcsr.scala 315:32:@2003.4]
  wire  mip_SSIP; // @[rvcsr.scala 315:32:@2005.4]
  wire  mip_rsrvd4; // @[rvcsr.scala 315:32:@2007.4]
  wire  _T_367; // @[rvcsr.scala 315:32:@2009.4]
  wire  mip_UTIP; // @[rvcsr.scala 315:32:@2011.4]
  wire  mip_STIP; // @[rvcsr.scala 315:32:@2013.4]
  wire  mip_rsrvd3; // @[rvcsr.scala 315:32:@2015.4]
  wire  _T_371; // @[rvcsr.scala 315:32:@2017.4]
  wire  mip_UEIP; // @[rvcsr.scala 315:32:@2019.4]
  wire  mip_SEIP; // @[rvcsr.scala 315:32:@2021.4]
  wire  mip_rsrvd2; // @[rvcsr.scala 315:32:@2023.4]
  wire  mip_MEIP; // @[rvcsr.scala 315:32:@2025.4]
  wire [18:0] mip_rsrvd1; // @[rvcsr.scala 315:32:@2027.4]
  wire [1:0] _T_383; // @[rvcsr.scala 317:34:@2046.4]
  wire  _T_384; // @[rvcsr.scala 317:34:@2048.4]
  wire [2:0] _T_385; // @[rvcsr.scala 317:34:@2050.4]
  wire [2:0] _T_386; // @[rvcsr.scala 317:34:@2052.4]
  wire  _T_387; // @[rvcsr.scala 317:34:@2054.4]
  wire  _T_388; // @[rvcsr.scala 317:34:@2056.4]
  wire  _T_389; // @[rvcsr.scala 317:34:@2058.4]
  wire  _T_390; // @[rvcsr.scala 317:34:@2060.4]
  wire  _T_391; // @[rvcsr.scala 317:34:@2062.4]
  wire  _T_392; // @[rvcsr.scala 317:34:@2064.4]
  wire  _T_393; // @[rvcsr.scala 317:34:@2066.4]
  wire [11:0] _T_394; // @[rvcsr.scala 317:34:@2068.4]
  wire [3:0] _T_395; // @[rvcsr.scala 317:34:@2070.4]
  wire [1:0] csr_priv; // @[rvcsr.scala 319:27:@2085.4]
  wire  legal_priv; // @[rvcsr.scala 320:28:@2086.4]
  wire  priv_inst; // @[rvcsr.scala 321:28:@2087.4]
  wire [2:0] priv_inst_type; // @[rvcsr.scala 322:33:@2088.4]
  wire  _T_396; // @[rvcsr.scala 323:33:@2089.4]
  wire  _T_398; // @[rvcsr.scala 323:61:@2090.4]
  wire  inst_ecall; // @[rvcsr.scala 323:44:@2091.4]
  wire  _T_401; // @[rvcsr.scala 324:62:@2093.4]
  wire  inst_ebreak; // @[rvcsr.scala 324:45:@2094.4]
  wire  _T_404; // @[rvcsr.scala 325:59:@2096.4]
  wire  inst_ret; // @[rvcsr.scala 325:42:@2097.4]
  wire  _T_405; // @[rvcsr.scala 328:31:@2098.4]
  wire  _T_406; // @[rvcsr.scala 328:45:@2099.4]
  wire  _T_407; // @[rvcsr.scala 331:21:@2101.4]
  wire [1:0] _T_409; // @[rvcsr.scala 333:24:@2104.6]
  wire [2:0] _T_410; // @[rvcsr.scala 333:24:@2105.6]
  wire [1:0] _T_411; // @[rvcsr.scala 333:24:@2106.6]
  wire  _T_690; // @[rvcsr.scala 382:28:@2294.4]
  wire  _T_691; // @[rvcsr.scala 382:40:@2295.4]
  wire  read_only; // @[rvcsr.scala 382:32:@2296.4]
  wire  _T_693; // @[rvcsr.scala 384:20:@2298.4]
  wire  _T_695; // @[rvcsr.scala 384:33:@2299.4]
  wire  _T_696; // @[rvcsr.scala 384:31:@2300.4]
  wire  csr_wen; // @[rvcsr.scala 384:43:@2301.4]
  wire  _T_491; // @[rvcsr.scala 380:61:@2194.4]
  wire  _T_1046; // @[rvcsr.scala 392:30:@2535.4]
  wire [31:0] _T_1048; // @[rvcsr.scala 392:22:@2536.4]
  wire  _T_1049; // @[rvcsr.scala 392:73:@2537.4]
  wire [31:0] _T_1051; // @[rvcsr.scala 392:65:@2538.4]
  wire [31:0] _T_1052; // @[rvcsr.scala 392:60:@2539.4]
  wire  _T_1053; // @[rvcsr.scala 392:119:@2540.4]
  wire [31:0] _T_1055; // @[rvcsr.scala 392:111:@2541.4]
  wire [31:0] _T_1056; // @[rvcsr.scala 392:107:@2542.4]
  wire [31:0] csr_wdata; // @[rvcsr.scala 392:104:@2543.4]
  wire [30:0] _T_1152; // @[:@2688.8]
  wire  _T_1156; // @[rvcsr.scala 435:47:@2696.8]
  wire  _GEN_67; // @[rvcsr.scala 434:37:@2686.6]
  wire  mip_MSIP; // @[rvcsr.scala 393:19:@2545.4]
  wire [2:0] _T_412; // @[rvcsr.scala 333:24:@2107.6]
  wire [5:0] _T_413; // @[rvcsr.scala 333:24:@2108.6]
  wire  _T_1160; // @[rvcsr.scala 435:47:@2704.8]
  wire  _GEN_32; // @[rvcsr.scala 331:38:@2102.4]
  wire  _GEN_66; // @[rvcsr.scala 434:37:@2686.6]
  wire  mip_MTIP; // @[rvcsr.scala 393:19:@2545.4]
  wire [1:0] _T_414; // @[rvcsr.scala 333:24:@2109.6]
  wire [2:0] _T_415; // @[rvcsr.scala 333:24:@2110.6]
  wire [1:0] _T_416; // @[rvcsr.scala 333:24:@2111.6]
  wire [19:0] _T_417; // @[rvcsr.scala 333:24:@2112.6]
  wire [21:0] _T_418; // @[rvcsr.scala 333:24:@2113.6]
  wire [24:0] _T_419; // @[rvcsr.scala 333:24:@2114.6]
  wire [30:0] _T_420; // @[rvcsr.scala 333:24:@2115.6]
  wire [31:0] _GEN_33; // @[rvcsr.scala 331:38:@2102.4]
  wire  _T_421; // @[rvcsr.scala 337:32:@2118.4]
  wire  _T_422; // @[rvcsr.scala 337:20:@2119.4]
  wire  _T_425; // @[rvcsr.scala 337:61:@2121.4]
  wire  _T_426; // @[rvcsr.scala 337:46:@2122.4]
  wire  mstatus_SIE; // @[rvcsr.scala 531:26:@3212.4]
  wire  mstatus_UIE; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _T_428; // @[rvcsr.scala 342:32:@2128.6]
  wire  mstatus_UPIE; // @[rvcsr.scala 531:26:@3212.4]
  wire  _T_469; // @[rvcsr.scala 380:61:@2183.4]
  wire  _T_1066; // @[rvcsr.scala 396:55:@2556.8]
  wire  _T_1070; // @[rvcsr.scala 396:55:@2564.8]
  wire  _GEN_35; // @[rvcsr.scala 337:73:@2123.4]
  wire  _GEN_55; // @[rvcsr.scala 395:41:@2546.6]
  wire  _GEN_173; // @[rvcsr.scala 393:19:@2545.4]
  wire  mstatus_MPIE; // @[rvcsr.scala 531:26:@3212.4]
  wire  _GEN_34; // @[rvcsr.scala 337:73:@2123.4]
  wire  _GEN_54; // @[rvcsr.scala 395:41:@2546.6]
  wire  _GEN_172; // @[rvcsr.scala 393:19:@2545.4]
  wire  mstatus_MIE; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _T_429; // @[rvcsr.scala 342:32:@2129.6]
  wire  mstatus_rsrvd4; // @[rvcsr.scala 531:26:@3212.4]
  wire [2:0] _T_430; // @[rvcsr.scala 342:32:@2130.6]
  wire [4:0] _T_431; // @[rvcsr.scala 342:32:@2131.6]
  wire  mstatus_rsrvd3; // @[rvcsr.scala 531:26:@3212.4]
  wire  mstatus_SPIE; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _T_432; // @[rvcsr.scala 342:32:@2132.6]
  wire [1:0] mstatus_rsrvd2; // @[rvcsr.scala 531:26:@3212.4]
  wire  mstatus_SPP; // @[rvcsr.scala 531:26:@3212.4]
  wire [2:0] _T_433; // @[rvcsr.scala 342:32:@2133.6]
  wire [3:0] _T_434; // @[rvcsr.scala 342:32:@2134.6]
  wire [5:0] _T_435; // @[rvcsr.scala 342:32:@2135.6]
  wire [10:0] _T_436; // @[rvcsr.scala 342:32:@2136.6]
  wire [1:0] mstatus_FS; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] mstatus_MPP; // @[rvcsr.scala 531:26:@3212.4]
  wire [3:0] _T_437; // @[rvcsr.scala 342:32:@2137.6]
  wire  mstatus_SUM; // @[rvcsr.scala 531:26:@3212.4]
  wire  mstatus_MPRV; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _T_438; // @[rvcsr.scala 342:32:@2138.6]
  wire [1:0] mstatus_XS; // @[rvcsr.scala 531:26:@3212.4]
  wire [3:0] _T_439; // @[rvcsr.scala 342:32:@2139.6]
  wire [7:0] _T_440; // @[rvcsr.scala 342:32:@2140.6]
  wire  mstatus_TW; // @[rvcsr.scala 531:26:@3212.4]
  wire  mstatus_TVM; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _T_441; // @[rvcsr.scala 342:32:@2141.6]
  wire  mstatus_MXR; // @[rvcsr.scala 531:26:@3212.4]
  wire [2:0] _T_442; // @[rvcsr.scala 342:32:@2142.6]
  wire  mstatus_SD; // @[rvcsr.scala 531:26:@3212.4]
  wire [7:0] mstatus_rsrvd1; // @[rvcsr.scala 531:26:@3212.4]
  wire [8:0] _T_443; // @[rvcsr.scala 342:32:@2143.6]
  wire  mstatus_TSR; // @[rvcsr.scala 531:26:@3212.4]
  wire [9:0] _T_444; // @[rvcsr.scala 342:32:@2144.6]
  wire [12:0] _T_445; // @[rvcsr.scala 342:32:@2145.6]
  wire [20:0] _T_446; // @[rvcsr.scala 342:32:@2146.6]
  wire [31:0] _T_447; // @[rvcsr.scala 342:32:@2147.6]
  wire [1:0] _GEN_36; // @[rvcsr.scala 337:73:@2123.4]
  wire [31:0] _GEN_38; // @[rvcsr.scala 337:73:@2123.4]
  wire [31:0] _GEN_39; // @[rvcsr.scala 346:21:@2150.4]
  wire [31:0] _GEN_40; // @[rvcsr.scala 346:21:@2150.4]
  wire  _T_509; // @[rvcsr.scala 380:61:@2203.4]
  wire  _T_1325; // @[rvcsr.scala 511:49:@3179.8]
  wire  _GEN_167; // @[rvcsr.scala 510:38:@3155.6]
  wire  _GEN_252; // @[rvcsr.scala 393:19:@2545.4]
  wire  dcsr_ebreakm; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_42; // @[rvcsr.scala 352:22:@2154.4]
  wire [31:0] _GEN_43; // @[rvcsr.scala 352:22:@2154.4]
  wire  _T_456; // @[rvcsr.scala 361:46:@2165.4]
  wire [1:0] dcsr_prv; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _GEN_46; // @[rvcsr.scala 361:72:@2166.4]
  wire [31:0] _GEN_47; // @[rvcsr.scala 361:72:@2166.4]
  wire  _T_458; // @[Conditional.scala 37:30:@2172.6]
  wire [31:0] _GEN_48; // @[Conditional.scala 40:58:@2173.6]
  wire [31:0] _GEN_49; // @[Conditional.scala 40:58:@2173.6]
  wire [31:0] _GEN_50; // @[Conditional.scala 40:58:@2173.6]
  wire [31:0] _GEN_51; // @[rvcsr.scala 368:25:@2171.4]
  wire [31:0] _GEN_52; // @[rvcsr.scala 368:25:@2171.4]
  wire [31:0] _GEN_53; // @[rvcsr.scala 368:25:@2171.4]
  wire  _T_473; // @[rvcsr.scala 380:61:@2185.4]
  wire  _T_475; // @[rvcsr.scala 380:61:@2186.4]
  wire  _T_477; // @[rvcsr.scala 380:61:@2187.4]
  wire  _T_479; // @[rvcsr.scala 380:61:@2188.4]
  wire  _T_481; // @[rvcsr.scala 380:61:@2189.4]
  wire  _T_483; // @[rvcsr.scala 380:61:@2190.4]
  wire  _T_485; // @[rvcsr.scala 380:61:@2191.4]
  wire  _T_487; // @[rvcsr.scala 380:61:@2192.4]
  wire  _T_489; // @[rvcsr.scala 380:61:@2193.4]
  wire  _T_493; // @[rvcsr.scala 380:61:@2195.4]
  wire  _T_495; // @[rvcsr.scala 380:61:@2196.4]
  wire  _T_497; // @[rvcsr.scala 380:61:@2197.4]
  wire  _T_499; // @[rvcsr.scala 380:61:@2198.4]
  wire  _T_501; // @[rvcsr.scala 380:61:@2199.4]
  wire  _T_503; // @[rvcsr.scala 380:61:@2200.4]
  wire  _T_505; // @[rvcsr.scala 380:61:@2201.4]
  wire  _T_507; // @[rvcsr.scala 380:61:@2202.4]
  wire  _T_511; // @[rvcsr.scala 380:61:@2204.4]
  wire  _T_513; // @[rvcsr.scala 380:61:@2205.4]
  wire  _T_515; // @[rvcsr.scala 380:61:@2206.4]
  wire  _T_517; // @[rvcsr.scala 380:61:@2207.4]
  wire  _T_519; // @[rvcsr.scala 380:61:@2208.4]
  wire  _T_521; // @[rvcsr.scala 380:61:@2209.4]
  wire  _T_523; // @[rvcsr.scala 380:61:@2210.4]
  wire  _T_525; // @[rvcsr.scala 380:61:@2211.4]
  wire  _T_527; // @[rvcsr.scala 380:61:@2212.4]
  wire  _T_529; // @[rvcsr.scala 380:61:@2213.4]
  wire  _T_531; // @[rvcsr.scala 380:61:@2214.4]
  wire  _T_533; // @[rvcsr.scala 380:61:@2215.4]
  wire  _T_535; // @[rvcsr.scala 380:61:@2216.4]
  wire  _T_537; // @[rvcsr.scala 380:61:@2217.4]
  wire  _T_539; // @[rvcsr.scala 380:61:@2218.4]
  wire  _T_541; // @[rvcsr.scala 380:61:@2219.4]
  wire  _T_543; // @[rvcsr.scala 380:61:@2220.4]
  wire  _T_545; // @[rvcsr.scala 380:61:@2221.4]
  wire  _T_547; // @[rvcsr.scala 380:61:@2222.4]
  wire  _T_549; // @[rvcsr.scala 380:61:@2223.4]
  wire  _T_551; // @[rvcsr.scala 380:61:@2224.4]
  wire  _T_553; // @[rvcsr.scala 380:61:@2225.4]
  wire  _T_555; // @[rvcsr.scala 380:61:@2226.4]
  wire  _T_557; // @[rvcsr.scala 380:61:@2227.4]
  wire  _T_559; // @[rvcsr.scala 380:61:@2228.4]
  wire  _T_561; // @[rvcsr.scala 380:61:@2229.4]
  wire  _T_563; // @[rvcsr.scala 380:61:@2230.4]
  wire  _T_565; // @[rvcsr.scala 380:61:@2231.4]
  wire  _T_567; // @[rvcsr.scala 380:61:@2232.4]
  wire  _T_569; // @[rvcsr.scala 380:61:@2233.4]
  wire  _T_571; // @[rvcsr.scala 380:61:@2234.4]
  wire  _T_573; // @[rvcsr.scala 380:61:@2235.4]
  wire  _T_575; // @[rvcsr.scala 380:61:@2236.4]
  wire  _T_577; // @[rvcsr.scala 380:61:@2237.4]
  wire  _T_579; // @[rvcsr.scala 380:61:@2238.4]
  wire  _T_581; // @[rvcsr.scala 380:61:@2239.4]
  wire  _T_583; // @[rvcsr.scala 380:61:@2240.4]
  wire  _T_585; // @[rvcsr.scala 380:61:@2241.4]
  wire  _T_587; // @[rvcsr.scala 380:61:@2242.4]
  wire  _T_589; // @[rvcsr.scala 380:61:@2243.4]
  wire  _T_591; // @[rvcsr.scala 380:61:@2244.4]
  wire  _T_593; // @[rvcsr.scala 380:61:@2245.4]
  wire  _T_595; // @[rvcsr.scala 380:61:@2246.4]
  wire  _T_597; // @[rvcsr.scala 380:61:@2247.4]
  wire  _T_599; // @[rvcsr.scala 380:61:@2248.4]
  wire  _T_601; // @[rvcsr.scala 380:61:@2249.4]
  wire  _T_603; // @[rvcsr.scala 380:61:@2250.4]
  wire  _T_605; // @[rvcsr.scala 380:61:@2251.4]
  wire  _T_607; // @[rvcsr.scala 380:61:@2252.4]
  wire  _T_609; // @[rvcsr.scala 380:61:@2253.4]
  wire  _T_611; // @[rvcsr.scala 380:61:@2254.4]
  wire  _T_613; // @[rvcsr.scala 380:61:@2255.4]
  wire  _T_615; // @[rvcsr.scala 380:61:@2256.4]
  wire  _T_617; // @[rvcsr.scala 380:61:@2257.4]
  wire  _T_619; // @[rvcsr.scala 380:61:@2258.4]
  wire  _T_621; // @[rvcsr.scala 380:61:@2259.4]
  wire  _T_623; // @[rvcsr.scala 380:61:@2260.4]
  wire  _T_625; // @[rvcsr.scala 380:61:@2261.4]
  wire  _T_627; // @[rvcsr.scala 380:61:@2262.4]
  wire  _T_629; // @[rvcsr.scala 380:61:@2263.4]
  wire  _T_631; // @[rvcsr.scala 380:61:@2264.4]
  wire  _T_633; // @[rvcsr.scala 380:61:@2265.4]
  wire  _T_635; // @[rvcsr.scala 380:61:@2266.4]
  wire  _T_637; // @[rvcsr.scala 380:61:@2267.4]
  wire  _T_639; // @[rvcsr.scala 380:61:@2268.4]
  wire  _T_641; // @[rvcsr.scala 380:61:@2269.4]
  wire  _T_643; // @[rvcsr.scala 380:61:@2270.4]
  wire  _T_645; // @[rvcsr.scala 380:61:@2271.4]
  wire  _T_647; // @[rvcsr.scala 380:61:@2272.4]
  wire  _T_649; // @[rvcsr.scala 380:61:@2273.4]
  wire  _T_651; // @[rvcsr.scala 380:61:@2274.4]
  wire  _T_653; // @[rvcsr.scala 380:61:@2275.4]
  wire  _T_655; // @[rvcsr.scala 380:61:@2276.4]
  wire  _T_657; // @[rvcsr.scala 380:61:@2277.4]
  wire  _T_659; // @[rvcsr.scala 380:61:@2278.4]
  wire  _T_661; // @[rvcsr.scala 380:61:@2279.4]
  wire  _T_663; // @[rvcsr.scala 380:61:@2280.4]
  wire  _T_665; // @[rvcsr.scala 380:61:@2281.4]
  wire  _T_667; // @[rvcsr.scala 380:61:@2282.4]
  wire  _T_669; // @[rvcsr.scala 380:61:@2283.4]
  wire  _T_671; // @[rvcsr.scala 380:61:@2284.4]
  wire  _T_673; // @[rvcsr.scala 380:61:@2285.4]
  wire  _T_675; // @[rvcsr.scala 380:61:@2286.4]
  wire  _T_677; // @[rvcsr.scala 380:61:@2287.4]
  wire  _T_679; // @[rvcsr.scala 380:61:@2288.4]
  wire  _T_681; // @[rvcsr.scala 380:61:@2289.4]
  wire  _T_683; // @[rvcsr.scala 380:61:@2290.4]
  wire  _T_685; // @[rvcsr.scala 380:61:@2291.4]
  wire  _T_687; // @[rvcsr.scala 380:61:@2292.4]
  wire  _T_689; // @[rvcsr.scala 380:61:@2293.4]
  wire  _T_813; // @[Mux.scala 46:19:@2302.4]
  wire [31:0] _T_814; // @[Mux.scala 46:16:@2303.4]
  wire  _T_815; // @[Mux.scala 46:19:@2304.4]
  wire [31:0] _T_816; // @[Mux.scala 46:16:@2305.4]
  wire  _T_817; // @[Mux.scala 46:19:@2306.4]
  wire [31:0] _T_818; // @[Mux.scala 46:16:@2307.4]
  wire  _T_819; // @[Mux.scala 46:19:@2308.4]
  wire [31:0] _T_820; // @[Mux.scala 46:16:@2309.4]
  wire  _T_821; // @[Mux.scala 46:19:@2310.4]
  wire [31:0] _T_822; // @[Mux.scala 46:16:@2311.4]
  wire  _T_823; // @[Mux.scala 46:19:@2312.4]
  wire [31:0] _T_824; // @[Mux.scala 46:16:@2313.4]
  wire  _T_825; // @[Mux.scala 46:19:@2314.4]
  wire [31:0] _T_826; // @[Mux.scala 46:16:@2315.4]
  wire  _T_827; // @[Mux.scala 46:19:@2316.4]
  wire [31:0] _T_828; // @[Mux.scala 46:16:@2317.4]
  wire  _T_829; // @[Mux.scala 46:19:@2318.4]
  wire [31:0] _T_830; // @[Mux.scala 46:16:@2319.4]
  wire  _T_831; // @[Mux.scala 46:19:@2320.4]
  wire [31:0] _T_832; // @[Mux.scala 46:16:@2321.4]
  wire  _T_833; // @[Mux.scala 46:19:@2322.4]
  wire [31:0] _T_834; // @[Mux.scala 46:16:@2323.4]
  wire  _T_835; // @[Mux.scala 46:19:@2324.4]
  wire [31:0] _T_836; // @[Mux.scala 46:16:@2325.4]
  wire  _T_837; // @[Mux.scala 46:19:@2326.4]
  wire [31:0] _T_838; // @[Mux.scala 46:16:@2327.4]
  wire  _T_839; // @[Mux.scala 46:19:@2328.4]
  wire [31:0] _T_840; // @[Mux.scala 46:16:@2329.4]
  wire  _T_841; // @[Mux.scala 46:19:@2330.4]
  wire [31:0] _T_842; // @[Mux.scala 46:16:@2331.4]
  wire  _T_843; // @[Mux.scala 46:19:@2332.4]
  wire [31:0] _T_844; // @[Mux.scala 46:16:@2333.4]
  wire  _T_845; // @[Mux.scala 46:19:@2334.4]
  wire [31:0] _T_846; // @[Mux.scala 46:16:@2335.4]
  wire  _T_847; // @[Mux.scala 46:19:@2336.4]
  wire [31:0] _T_848; // @[Mux.scala 46:16:@2337.4]
  wire  _T_849; // @[Mux.scala 46:19:@2338.4]
  wire [31:0] _T_850; // @[Mux.scala 46:16:@2339.4]
  wire  _T_851; // @[Mux.scala 46:19:@2340.4]
  wire [31:0] _T_852; // @[Mux.scala 46:16:@2341.4]
  wire  _T_853; // @[Mux.scala 46:19:@2342.4]
  wire [31:0] _T_854; // @[Mux.scala 46:16:@2343.4]
  wire  _T_855; // @[Mux.scala 46:19:@2344.4]
  wire [31:0] _T_856; // @[Mux.scala 46:16:@2345.4]
  wire  _T_857; // @[Mux.scala 46:19:@2346.4]
  wire [31:0] _T_858; // @[Mux.scala 46:16:@2347.4]
  wire  _T_859; // @[Mux.scala 46:19:@2348.4]
  wire [31:0] _T_860; // @[Mux.scala 46:16:@2349.4]
  wire  _T_861; // @[Mux.scala 46:19:@2350.4]
  wire [31:0] _T_862; // @[Mux.scala 46:16:@2351.4]
  wire  _T_863; // @[Mux.scala 46:19:@2352.4]
  wire [31:0] _T_864; // @[Mux.scala 46:16:@2353.4]
  wire  _T_865; // @[Mux.scala 46:19:@2354.4]
  wire [31:0] _T_866; // @[Mux.scala 46:16:@2355.4]
  wire  _T_867; // @[Mux.scala 46:19:@2356.4]
  wire [31:0] _T_868; // @[Mux.scala 46:16:@2357.4]
  wire  _T_869; // @[Mux.scala 46:19:@2358.4]
  wire [31:0] _T_870; // @[Mux.scala 46:16:@2359.4]
  wire  _T_871; // @[Mux.scala 46:19:@2360.4]
  wire [31:0] _T_872; // @[Mux.scala 46:16:@2361.4]
  wire  _T_873; // @[Mux.scala 46:19:@2362.4]
  wire [31:0] _T_874; // @[Mux.scala 46:16:@2363.4]
  wire  _T_875; // @[Mux.scala 46:19:@2364.4]
  wire [31:0] _T_876; // @[Mux.scala 46:16:@2365.4]
  wire  _T_877; // @[Mux.scala 46:19:@2366.4]
  wire [31:0] _T_878; // @[Mux.scala 46:16:@2367.4]
  wire  _T_879; // @[Mux.scala 46:19:@2368.4]
  wire [31:0] _T_880; // @[Mux.scala 46:16:@2369.4]
  wire  _T_881; // @[Mux.scala 46:19:@2370.4]
  wire [31:0] _T_882; // @[Mux.scala 46:16:@2371.4]
  wire  _T_883; // @[Mux.scala 46:19:@2372.4]
  wire [31:0] _T_884; // @[Mux.scala 46:16:@2373.4]
  wire  _T_885; // @[Mux.scala 46:19:@2374.4]
  wire [31:0] _T_886; // @[Mux.scala 46:16:@2375.4]
  wire  _T_887; // @[Mux.scala 46:19:@2376.4]
  wire [31:0] _T_888; // @[Mux.scala 46:16:@2377.4]
  wire  _T_889; // @[Mux.scala 46:19:@2378.4]
  wire [31:0] _T_890; // @[Mux.scala 46:16:@2379.4]
  wire  _T_891; // @[Mux.scala 46:19:@2380.4]
  wire [31:0] _T_892; // @[Mux.scala 46:16:@2381.4]
  wire  _T_893; // @[Mux.scala 46:19:@2382.4]
  wire [31:0] _T_894; // @[Mux.scala 46:16:@2383.4]
  wire  _T_895; // @[Mux.scala 46:19:@2384.4]
  wire [31:0] _T_896; // @[Mux.scala 46:16:@2385.4]
  wire  _T_897; // @[Mux.scala 46:19:@2386.4]
  wire [31:0] _T_898; // @[Mux.scala 46:16:@2387.4]
  wire  _T_899; // @[Mux.scala 46:19:@2388.4]
  wire [31:0] _T_900; // @[Mux.scala 46:16:@2389.4]
  wire  _T_901; // @[Mux.scala 46:19:@2390.4]
  wire [31:0] _T_902; // @[Mux.scala 46:16:@2391.4]
  wire  _T_903; // @[Mux.scala 46:19:@2392.4]
  wire [31:0] _T_904; // @[Mux.scala 46:16:@2393.4]
  wire  _T_905; // @[Mux.scala 46:19:@2394.4]
  wire [31:0] _T_906; // @[Mux.scala 46:16:@2395.4]
  wire  _T_907; // @[Mux.scala 46:19:@2396.4]
  wire [31:0] _T_908; // @[Mux.scala 46:16:@2397.4]
  wire  _T_909; // @[Mux.scala 46:19:@2398.4]
  wire [31:0] _T_910; // @[Mux.scala 46:16:@2399.4]
  wire  _T_911; // @[Mux.scala 46:19:@2400.4]
  wire [31:0] _T_912; // @[Mux.scala 46:16:@2401.4]
  wire  _T_913; // @[Mux.scala 46:19:@2402.4]
  wire [31:0] _T_914; // @[Mux.scala 46:16:@2403.4]
  wire  _T_915; // @[Mux.scala 46:19:@2404.4]
  wire [31:0] _T_916; // @[Mux.scala 46:16:@2405.4]
  wire  _T_917; // @[Mux.scala 46:19:@2406.4]
  wire [31:0] _T_918; // @[Mux.scala 46:16:@2407.4]
  wire  _T_919; // @[Mux.scala 46:19:@2408.4]
  wire [31:0] _T_920; // @[Mux.scala 46:16:@2409.4]
  wire  _T_921; // @[Mux.scala 46:19:@2410.4]
  wire [31:0] _T_922; // @[Mux.scala 46:16:@2411.4]
  wire  _T_923; // @[Mux.scala 46:19:@2412.4]
  wire [31:0] _T_924; // @[Mux.scala 46:16:@2413.4]
  wire  _T_925; // @[Mux.scala 46:19:@2414.4]
  wire [31:0] _T_926; // @[Mux.scala 46:16:@2415.4]
  wire  _T_927; // @[Mux.scala 46:19:@2416.4]
  wire [31:0] _T_928; // @[Mux.scala 46:16:@2417.4]
  wire  _T_929; // @[Mux.scala 46:19:@2418.4]
  wire [31:0] _T_930; // @[Mux.scala 46:16:@2419.4]
  wire  _T_931; // @[Mux.scala 46:19:@2420.4]
  wire [31:0] _T_932; // @[Mux.scala 46:16:@2421.4]
  wire  _T_933; // @[Mux.scala 46:19:@2422.4]
  wire [31:0] _T_934; // @[Mux.scala 46:16:@2423.4]
  wire  _T_935; // @[Mux.scala 46:19:@2424.4]
  wire [31:0] _T_936; // @[Mux.scala 46:16:@2425.4]
  wire  _T_937; // @[Mux.scala 46:19:@2426.4]
  wire [31:0] _T_938; // @[Mux.scala 46:16:@2427.4]
  wire  _T_939; // @[Mux.scala 46:19:@2428.4]
  wire [31:0] _T_940; // @[Mux.scala 46:16:@2429.4]
  wire  _T_941; // @[Mux.scala 46:19:@2430.4]
  wire [31:0] _T_942; // @[Mux.scala 46:16:@2431.4]
  wire  _T_943; // @[Mux.scala 46:19:@2432.4]
  wire [31:0] _T_944; // @[Mux.scala 46:16:@2433.4]
  wire  _T_945; // @[Mux.scala 46:19:@2434.4]
  wire [31:0] _T_946; // @[Mux.scala 46:16:@2435.4]
  wire  _T_947; // @[Mux.scala 46:19:@2436.4]
  wire [31:0] _T_948; // @[Mux.scala 46:16:@2437.4]
  wire  _T_949; // @[Mux.scala 46:19:@2438.4]
  wire [31:0] _T_950; // @[Mux.scala 46:16:@2439.4]
  wire  _T_951; // @[Mux.scala 46:19:@2440.4]
  wire [31:0] _T_952; // @[Mux.scala 46:16:@2441.4]
  wire  _T_953; // @[Mux.scala 46:19:@2442.4]
  wire [31:0] _T_954; // @[Mux.scala 46:16:@2443.4]
  wire  _T_955; // @[Mux.scala 46:19:@2444.4]
  wire [31:0] _T_956; // @[Mux.scala 46:16:@2445.4]
  wire  _T_957; // @[Mux.scala 46:19:@2446.4]
  wire [31:0] _T_958; // @[Mux.scala 46:16:@2447.4]
  wire  _T_959; // @[Mux.scala 46:19:@2448.4]
  wire [31:0] _T_960; // @[Mux.scala 46:16:@2449.4]
  wire  _T_961; // @[Mux.scala 46:19:@2450.4]
  wire [31:0] _T_962; // @[Mux.scala 46:16:@2451.4]
  wire  _T_963; // @[Mux.scala 46:19:@2452.4]
  wire [31:0] _T_964; // @[Mux.scala 46:16:@2453.4]
  wire  _T_965; // @[Mux.scala 46:19:@2454.4]
  wire [31:0] _T_966; // @[Mux.scala 46:16:@2455.4]
  wire  _T_967; // @[Mux.scala 46:19:@2456.4]
  wire [31:0] _T_968; // @[Mux.scala 46:16:@2457.4]
  wire  _T_969; // @[Mux.scala 46:19:@2458.4]
  wire [31:0] _T_970; // @[Mux.scala 46:16:@2459.4]
  wire  _T_971; // @[Mux.scala 46:19:@2460.4]
  wire [31:0] _T_972; // @[Mux.scala 46:16:@2461.4]
  wire  _T_973; // @[Mux.scala 46:19:@2462.4]
  wire [31:0] _T_974; // @[Mux.scala 46:16:@2463.4]
  wire  _T_975; // @[Mux.scala 46:19:@2464.4]
  wire [31:0] _T_976; // @[Mux.scala 46:16:@2465.4]
  wire  _T_977; // @[Mux.scala 46:19:@2466.4]
  wire [31:0] _T_978; // @[Mux.scala 46:16:@2467.4]
  wire  _T_979; // @[Mux.scala 46:19:@2468.4]
  wire [31:0] _T_980; // @[Mux.scala 46:16:@2469.4]
  wire  _T_981; // @[Mux.scala 46:19:@2470.4]
  wire [31:0] _T_982; // @[Mux.scala 46:16:@2471.4]
  wire  _T_983; // @[Mux.scala 46:19:@2472.4]
  wire [31:0] _T_984; // @[Mux.scala 46:16:@2473.4]
  wire  _T_985; // @[Mux.scala 46:19:@2474.4]
  wire [31:0] _T_986; // @[Mux.scala 46:16:@2475.4]
  wire  _T_987; // @[Mux.scala 46:19:@2476.4]
  wire [31:0] _T_988; // @[Mux.scala 46:16:@2477.4]
  wire  _T_989; // @[Mux.scala 46:19:@2478.4]
  wire [31:0] _T_990; // @[Mux.scala 46:16:@2479.4]
  wire  _T_991; // @[Mux.scala 46:19:@2480.4]
  wire [31:0] _T_992; // @[Mux.scala 46:16:@2481.4]
  wire  _T_993; // @[Mux.scala 46:19:@2482.4]
  wire [31:0] _T_994; // @[Mux.scala 46:16:@2483.4]
  wire  _T_995; // @[Mux.scala 46:19:@2484.4]
  wire [31:0] _T_996; // @[Mux.scala 46:16:@2485.4]
  wire  _T_997; // @[Mux.scala 46:19:@2486.4]
  wire [31:0] _T_998; // @[Mux.scala 46:16:@2487.4]
  wire  _T_999; // @[Mux.scala 46:19:@2488.4]
  wire [31:0] _T_1000; // @[Mux.scala 46:16:@2489.4]
  wire  _T_1001; // @[Mux.scala 46:19:@2490.4]
  wire [31:0] _T_1002; // @[Mux.scala 46:16:@2491.4]
  wire  _T_1003; // @[Mux.scala 46:19:@2492.4]
  wire [31:0] _T_1004; // @[Mux.scala 46:16:@2493.4]
  wire  _T_1005; // @[Mux.scala 46:19:@2494.4]
  wire [31:0] _T_1006; // @[Mux.scala 46:16:@2495.4]
  wire  _T_1007; // @[Mux.scala 46:19:@2496.4]
  wire [31:0] _T_1008; // @[Mux.scala 46:16:@2497.4]
  wire  _T_1009; // @[Mux.scala 46:19:@2498.4]
  wire [31:0] _T_1010; // @[Mux.scala 46:16:@2499.4]
  wire  _T_1011; // @[Mux.scala 46:19:@2500.4]
  wire [31:0] _T_1012; // @[Mux.scala 46:16:@2501.4]
  wire  _T_1013; // @[Mux.scala 46:19:@2502.4]
  wire [31:0] _T_1014; // @[Mux.scala 46:16:@2503.4]
  wire  _T_1015; // @[Mux.scala 46:19:@2504.4]
  wire [31:0] _T_1016; // @[Mux.scala 46:16:@2505.4]
  wire  _T_1017; // @[Mux.scala 46:19:@2506.4]
  wire [31:0] _T_1018; // @[Mux.scala 46:16:@2507.4]
  wire  _T_1019; // @[Mux.scala 46:19:@2508.4]
  wire [31:0] _T_1020; // @[Mux.scala 46:16:@2509.4]
  wire  _T_1021; // @[Mux.scala 46:19:@2510.4]
  wire [31:0] _T_1022; // @[Mux.scala 46:16:@2511.4]
  wire  _T_1023; // @[Mux.scala 46:19:@2512.4]
  wire [31:0] _T_1024; // @[Mux.scala 46:16:@2513.4]
  wire  _T_1025; // @[Mux.scala 46:19:@2514.4]
  wire [31:0] _T_1026; // @[Mux.scala 46:16:@2515.4]
  wire  _T_1027; // @[Mux.scala 46:19:@2516.4]
  wire [31:0] _T_1028; // @[Mux.scala 46:16:@2517.4]
  wire  _T_1029; // @[Mux.scala 46:19:@2518.4]
  wire [31:0] _T_1030; // @[Mux.scala 46:16:@2519.4]
  wire  _T_1031; // @[Mux.scala 46:19:@2520.4]
  wire [31:0] _T_1032; // @[Mux.scala 46:16:@2521.4]
  wire  _T_1033; // @[Mux.scala 46:19:@2522.4]
  wire [31:0] _T_1034; // @[Mux.scala 46:16:@2523.4]
  wire  _T_1035; // @[Mux.scala 46:19:@2524.4]
  wire [31:0] _T_1036; // @[Mux.scala 46:16:@2525.4]
  wire  _T_1037; // @[Mux.scala 46:19:@2526.4]
  wire [31:0] _T_1038; // @[Mux.scala 46:16:@2527.4]
  wire  _T_1039; // @[Mux.scala 46:19:@2528.4]
  wire [31:0] _T_1040; // @[Mux.scala 46:16:@2529.4]
  wire  _T_1041; // @[Mux.scala 46:19:@2530.4]
  wire [31:0] _T_1042; // @[Mux.scala 46:16:@2531.4]
  wire [31:0] _T_1044; // @[rvcsr.scala 389:20:@2532.4]
  wire  _T_1065; // @[rvcsr.scala 396:55:@2554.8]
  wire [31:0] _GEN_56; // @[rvcsr.scala 395:41:@2546.6]
  wire [1:0] _T_1122; // @[rvcsr.scala 407:28:@2648.8]
  wire [2:0] _T_1123; // @[rvcsr.scala 407:28:@2649.8]
  wire [1:0] _T_1124; // @[rvcsr.scala 407:28:@2650.8]
  wire  _GEN_58; // @[rvcsr.scala 402:37:@2616.6]
  wire  mie_MSIE; // @[rvcsr.scala 393:19:@2545.4]
  wire [2:0] _T_1125; // @[rvcsr.scala 407:28:@2651.8]
  wire [5:0] _T_1126; // @[rvcsr.scala 407:28:@2652.8]
  wire  _GEN_57; // @[rvcsr.scala 402:37:@2616.6]
  wire  mie_MTIE; // @[rvcsr.scala 393:19:@2545.4]
  wire [1:0] _T_1127; // @[rvcsr.scala 407:28:@2653.8]
  wire [2:0] _T_1128; // @[rvcsr.scala 407:28:@2654.8]
  wire [1:0] _T_1129; // @[rvcsr.scala 407:28:@2655.8]
  wire [19:0] _T_1130; // @[rvcsr.scala 407:28:@2656.8]
  wire [21:0] _T_1131; // @[rvcsr.scala 407:28:@2657.8]
  wire [24:0] _T_1132; // @[rvcsr.scala 407:28:@2658.8]
  wire [30:0] _T_1133; // @[rvcsr.scala 407:28:@2659.8]
  wire [31:0] _GEN_59; // @[rvcsr.scala 402:37:@2616.6]
  wire [29:0] _T_1134; // @[rvcsr.scala 411:39:@2663.8]
  wire [31:0] _T_1140; // @[Cat.scala 30:58:@2665.8]
  wire [31:0] _GEN_60; // @[rvcsr.scala 410:39:@2662.6]
  wire [31:0] _GEN_61; // @[rvcsr.scala 414:44:@2668.6]
  wire [31:0] _GEN_62; // @[rvcsr.scala 418:42:@2671.6]
  wire [31:0] _GEN_63; // @[rvcsr.scala 422:38:@2674.6]
  wire [31:0] _GEN_64; // @[rvcsr.scala 426:40:@2680.6]
  wire [31:0] _GEN_65; // @[rvcsr.scala 430:39:@2683.6]
  wire [31:0] _GEN_68; // @[rvcsr.scala 434:37:@2686.6]
  wire [31:0] _T_1178; // @[rvcsr.scala 444:41:@2733.8]
  wire [63:0] _T_1179; // @[Cat.scala 30:58:@2734.8]
  wire [63:0] _GEN_69; // @[rvcsr.scala 442:40:@2732.6]
  wire [63:0] _T_1181; // @[Cat.scala 30:58:@2739.8]
  wire [63:0] _GEN_70; // @[rvcsr.scala 447:42:@2737.6]
  wire [63:0] _T_1183; // @[Cat.scala 30:58:@2744.8]
  wire [63:0] _GEN_71; // @[rvcsr.scala 452:41:@2742.6]
  wire [31:0] _T_1184; // @[rvcsr.scala 459:56:@2748.8]
  wire [63:0] _T_1185; // @[Cat.scala 30:58:@2749.8]
  wire [63:0] _GEN_72; // @[rvcsr.scala 457:43:@2747.6]
  wire [63:0] _T_1187; // @[Cat.scala 30:58:@2754.8]
  wire [63:0] _GEN_73; // @[rvcsr.scala 463:57:@2752.6]
  wire [63:0] _T_1189; // @[Cat.scala 30:58:@2759.8]
  wire [63:0] _GEN_74; // @[rvcsr.scala 463:57:@2757.6]
  wire [63:0] _T_1191; // @[Cat.scala 30:58:@2764.8]
  wire [63:0] _GEN_75; // @[rvcsr.scala 463:57:@2762.6]
  wire [63:0] _T_1193; // @[Cat.scala 30:58:@2769.8]
  wire [63:0] _GEN_76; // @[rvcsr.scala 463:57:@2767.6]
  wire [63:0] _T_1195; // @[Cat.scala 30:58:@2774.8]
  wire [63:0] _GEN_77; // @[rvcsr.scala 463:57:@2772.6]
  wire [63:0] _T_1197; // @[Cat.scala 30:58:@2779.8]
  wire [63:0] _GEN_78; // @[rvcsr.scala 463:57:@2777.6]
  wire [63:0] _T_1199; // @[Cat.scala 30:58:@2784.8]
  wire [63:0] _GEN_79; // @[rvcsr.scala 463:57:@2782.6]
  wire [63:0] _T_1201; // @[Cat.scala 30:58:@2789.8]
  wire [63:0] _GEN_80; // @[rvcsr.scala 463:57:@2787.6]
  wire [63:0] _T_1203; // @[Cat.scala 30:58:@2794.8]
  wire [63:0] _GEN_81; // @[rvcsr.scala 463:57:@2792.6]
  wire [63:0] _T_1205; // @[Cat.scala 30:58:@2799.8]
  wire [63:0] _GEN_82; // @[rvcsr.scala 463:57:@2797.6]
  wire [63:0] _T_1207; // @[Cat.scala 30:58:@2804.8]
  wire [63:0] _GEN_83; // @[rvcsr.scala 463:57:@2802.6]
  wire [63:0] _T_1209; // @[Cat.scala 30:58:@2809.8]
  wire [63:0] _GEN_84; // @[rvcsr.scala 463:57:@2807.6]
  wire [63:0] _T_1211; // @[Cat.scala 30:58:@2814.8]
  wire [63:0] _GEN_85; // @[rvcsr.scala 463:57:@2812.6]
  wire [63:0] _T_1213; // @[Cat.scala 30:58:@2819.8]
  wire [63:0] _GEN_86; // @[rvcsr.scala 463:57:@2817.6]
  wire [63:0] _T_1215; // @[Cat.scala 30:58:@2824.8]
  wire [63:0] _GEN_87; // @[rvcsr.scala 463:57:@2822.6]
  wire [63:0] _T_1217; // @[Cat.scala 30:58:@2829.8]
  wire [63:0] _GEN_88; // @[rvcsr.scala 463:57:@2827.6]
  wire [63:0] _T_1219; // @[Cat.scala 30:58:@2834.8]
  wire [63:0] _GEN_89; // @[rvcsr.scala 463:57:@2832.6]
  wire [63:0] _T_1221; // @[Cat.scala 30:58:@2839.8]
  wire [63:0] _GEN_90; // @[rvcsr.scala 463:57:@2837.6]
  wire [63:0] _T_1223; // @[Cat.scala 30:58:@2844.8]
  wire [63:0] _GEN_91; // @[rvcsr.scala 463:57:@2842.6]
  wire [63:0] _T_1225; // @[Cat.scala 30:58:@2849.8]
  wire [63:0] _GEN_92; // @[rvcsr.scala 463:57:@2847.6]
  wire [63:0] _T_1227; // @[Cat.scala 30:58:@2854.8]
  wire [63:0] _GEN_93; // @[rvcsr.scala 463:57:@2852.6]
  wire [63:0] _T_1229; // @[Cat.scala 30:58:@2859.8]
  wire [63:0] _GEN_94; // @[rvcsr.scala 463:57:@2857.6]
  wire [63:0] _T_1231; // @[Cat.scala 30:58:@2864.8]
  wire [63:0] _GEN_95; // @[rvcsr.scala 463:57:@2862.6]
  wire [63:0] _T_1233; // @[Cat.scala 30:58:@2869.8]
  wire [63:0] _GEN_96; // @[rvcsr.scala 463:57:@2867.6]
  wire [63:0] _T_1235; // @[Cat.scala 30:58:@2874.8]
  wire [63:0] _GEN_97; // @[rvcsr.scala 463:57:@2872.6]
  wire [63:0] _T_1237; // @[Cat.scala 30:58:@2879.8]
  wire [63:0] _GEN_98; // @[rvcsr.scala 463:57:@2877.6]
  wire [63:0] _T_1239; // @[Cat.scala 30:58:@2884.8]
  wire [63:0] _GEN_99; // @[rvcsr.scala 463:57:@2882.6]
  wire [63:0] _T_1241; // @[Cat.scala 30:58:@2889.8]
  wire [63:0] _GEN_100; // @[rvcsr.scala 463:57:@2887.6]
  wire [63:0] _T_1243; // @[Cat.scala 30:58:@2894.8]
  wire [63:0] _GEN_101; // @[rvcsr.scala 463:57:@2892.6]
  wire [63:0] _T_1245; // @[Cat.scala 30:58:@2899.8]
  wire [63:0] _GEN_102; // @[rvcsr.scala 470:58:@2897.6]
  wire [63:0] _T_1247; // @[Cat.scala 30:58:@2904.8]
  wire [63:0] _GEN_103; // @[rvcsr.scala 470:58:@2902.6]
  wire [63:0] _T_1249; // @[Cat.scala 30:58:@2909.8]
  wire [63:0] _GEN_104; // @[rvcsr.scala 470:58:@2907.6]
  wire [63:0] _T_1251; // @[Cat.scala 30:58:@2914.8]
  wire [63:0] _GEN_105; // @[rvcsr.scala 470:58:@2912.6]
  wire [63:0] _T_1253; // @[Cat.scala 30:58:@2919.8]
  wire [63:0] _GEN_106; // @[rvcsr.scala 470:58:@2917.6]
  wire [63:0] _T_1255; // @[Cat.scala 30:58:@2924.8]
  wire [63:0] _GEN_107; // @[rvcsr.scala 470:58:@2922.6]
  wire [63:0] _T_1257; // @[Cat.scala 30:58:@2929.8]
  wire [63:0] _GEN_108; // @[rvcsr.scala 470:58:@2927.6]
  wire [63:0] _T_1259; // @[Cat.scala 30:58:@2934.8]
  wire [63:0] _GEN_109; // @[rvcsr.scala 470:58:@2932.6]
  wire [63:0] _T_1261; // @[Cat.scala 30:58:@2939.8]
  wire [63:0] _GEN_110; // @[rvcsr.scala 470:58:@2937.6]
  wire [63:0] _T_1263; // @[Cat.scala 30:58:@2944.8]
  wire [63:0] _GEN_111; // @[rvcsr.scala 470:58:@2942.6]
  wire [63:0] _T_1265; // @[Cat.scala 30:58:@2949.8]
  wire [63:0] _GEN_112; // @[rvcsr.scala 470:58:@2947.6]
  wire [63:0] _T_1267; // @[Cat.scala 30:58:@2954.8]
  wire [63:0] _GEN_113; // @[rvcsr.scala 470:58:@2952.6]
  wire [63:0] _T_1269; // @[Cat.scala 30:58:@2959.8]
  wire [63:0] _GEN_114; // @[rvcsr.scala 470:58:@2957.6]
  wire [63:0] _T_1271; // @[Cat.scala 30:58:@2964.8]
  wire [63:0] _GEN_115; // @[rvcsr.scala 470:58:@2962.6]
  wire [63:0] _T_1273; // @[Cat.scala 30:58:@2969.8]
  wire [63:0] _GEN_116; // @[rvcsr.scala 470:58:@2967.6]
  wire [63:0] _T_1275; // @[Cat.scala 30:58:@2974.8]
  wire [63:0] _GEN_117; // @[rvcsr.scala 470:58:@2972.6]
  wire [63:0] _T_1277; // @[Cat.scala 30:58:@2979.8]
  wire [63:0] _GEN_118; // @[rvcsr.scala 470:58:@2977.6]
  wire [63:0] _T_1279; // @[Cat.scala 30:58:@2984.8]
  wire [63:0] _GEN_119; // @[rvcsr.scala 470:58:@2982.6]
  wire [63:0] _T_1281; // @[Cat.scala 30:58:@2989.8]
  wire [63:0] _GEN_120; // @[rvcsr.scala 470:58:@2987.6]
  wire [63:0] _T_1283; // @[Cat.scala 30:58:@2994.8]
  wire [63:0] _GEN_121; // @[rvcsr.scala 470:58:@2992.6]
  wire [63:0] _T_1285; // @[Cat.scala 30:58:@2999.8]
  wire [63:0] _GEN_122; // @[rvcsr.scala 470:58:@2997.6]
  wire [63:0] _T_1287; // @[Cat.scala 30:58:@3004.8]
  wire [63:0] _GEN_123; // @[rvcsr.scala 470:58:@3002.6]
  wire [63:0] _T_1289; // @[Cat.scala 30:58:@3009.8]
  wire [63:0] _GEN_124; // @[rvcsr.scala 470:58:@3007.6]
  wire [63:0] _T_1291; // @[Cat.scala 30:58:@3014.8]
  wire [63:0] _GEN_125; // @[rvcsr.scala 470:58:@3012.6]
  wire [63:0] _T_1293; // @[Cat.scala 30:58:@3019.8]
  wire [63:0] _GEN_126; // @[rvcsr.scala 470:58:@3017.6]
  wire [63:0] _T_1295; // @[Cat.scala 30:58:@3024.8]
  wire [63:0] _GEN_127; // @[rvcsr.scala 470:58:@3022.6]
  wire [63:0] _T_1297; // @[Cat.scala 30:58:@3029.8]
  wire [63:0] _GEN_128; // @[rvcsr.scala 470:58:@3027.6]
  wire [63:0] _T_1299; // @[Cat.scala 30:58:@3034.8]
  wire [63:0] _GEN_129; // @[rvcsr.scala 470:58:@3032.6]
  wire [63:0] _T_1301; // @[Cat.scala 30:58:@3039.8]
  wire [63:0] _GEN_130; // @[rvcsr.scala 470:58:@3037.6]
  wire [31:0] _GEN_131; // @[rvcsr.scala 477:55:@3042.6]
  wire [31:0] _GEN_132; // @[rvcsr.scala 477:55:@3045.6]
  wire [31:0] _GEN_133; // @[rvcsr.scala 477:55:@3048.6]
  wire [31:0] _GEN_134; // @[rvcsr.scala 477:55:@3051.6]
  wire [31:0] _GEN_135; // @[rvcsr.scala 477:55:@3054.6]
  wire [31:0] _GEN_136; // @[rvcsr.scala 477:55:@3057.6]
  wire [31:0] _GEN_137; // @[rvcsr.scala 477:55:@3060.6]
  wire [31:0] _GEN_138; // @[rvcsr.scala 477:55:@3063.6]
  wire [31:0] _GEN_139; // @[rvcsr.scala 477:55:@3066.6]
  wire [31:0] _GEN_140; // @[rvcsr.scala 477:55:@3069.6]
  wire [31:0] _GEN_141; // @[rvcsr.scala 477:55:@3072.6]
  wire [31:0] _GEN_142; // @[rvcsr.scala 477:55:@3075.6]
  wire [31:0] _GEN_143; // @[rvcsr.scala 477:55:@3078.6]
  wire [31:0] _GEN_144; // @[rvcsr.scala 477:55:@3081.6]
  wire [31:0] _GEN_145; // @[rvcsr.scala 477:55:@3084.6]
  wire [31:0] _GEN_146; // @[rvcsr.scala 477:55:@3087.6]
  wire [31:0] _GEN_147; // @[rvcsr.scala 477:55:@3090.6]
  wire [31:0] _GEN_148; // @[rvcsr.scala 477:55:@3093.6]
  wire [31:0] _GEN_149; // @[rvcsr.scala 477:55:@3096.6]
  wire [31:0] _GEN_150; // @[rvcsr.scala 477:55:@3099.6]
  wire [31:0] _GEN_151; // @[rvcsr.scala 477:55:@3102.6]
  wire [31:0] _GEN_152; // @[rvcsr.scala 477:55:@3105.6]
  wire [31:0] _GEN_153; // @[rvcsr.scala 477:55:@3108.6]
  wire [31:0] _GEN_154; // @[rvcsr.scala 477:55:@3111.6]
  wire [31:0] _GEN_155; // @[rvcsr.scala 477:55:@3114.6]
  wire [31:0] _GEN_156; // @[rvcsr.scala 477:55:@3117.6]
  wire [31:0] _GEN_157; // @[rvcsr.scala 477:55:@3120.6]
  wire [31:0] _GEN_158; // @[rvcsr.scala 477:55:@3123.6]
  wire [31:0] _GEN_159; // @[rvcsr.scala 477:55:@3126.6]
  wire [63:0] _T_1303; // @[Cat.scala 30:58:@3131.8]
  wire [63:0] _GEN_160; // @[rvcsr.scala 482:39:@3129.6]
  wire [63:0] _T_1305; // @[Cat.scala 30:58:@3136.8]
  wire [63:0] _GEN_161; // @[rvcsr.scala 487:42:@3134.6]
  wire [63:0] _T_1307; // @[Cat.scala 30:58:@3141.8]
  wire [63:0] _GEN_162; // @[rvcsr.scala 492:40:@3139.6]
  wire [31:0] _T_1308; // @[rvcsr.scala 499:56:@3145.8]
  wire [63:0] _T_1309; // @[Cat.scala 30:58:@3146.8]
  wire [63:0] _GEN_163; // @[rvcsr.scala 497:43:@3144.6]
  wire [31:0] _GEN_164; // @[rvcsr.scala 502:41:@3149.6]
  wire [31:0] _GEN_165; // @[rvcsr.scala 506:41:@3152.6]
  wire [2:0] dcsr_rsrvd3; // @[rvcsr.scala 531:26:@3212.4]
  wire  _GEN_166; // @[rvcsr.scala 510:38:@3155.6]
  wire  _GEN_251; // @[rvcsr.scala 393:19:@2545.4]
  wire  dcsr_step; // @[rvcsr.scala 531:26:@3212.4]
  wire [3:0] _T_1328; // @[rvcsr.scala 514:30:@3187.8]
  wire [5:0] _T_1329; // @[rvcsr.scala 514:30:@3188.8]
  wire  dcsr_stopcount; // @[rvcsr.scala 531:26:@3212.4]
  wire  dcsr_stoptime; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _T_1330; // @[rvcsr.scala 514:30:@3189.8]
  wire [2:0] dcsr_cause; // @[rvcsr.scala 531:26:@3212.4]
  wire [4:0] _T_1331; // @[rvcsr.scala 514:30:@3190.8]
  wire [10:0] _T_1332; // @[rvcsr.scala 514:30:@3191.8]
  wire  dcsr_ebreaks; // @[rvcsr.scala 531:26:@3212.4]
  wire  dcsr_ebreaku; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _T_1333; // @[rvcsr.scala 514:30:@3192.8]
  wire  dcsr_rsrvd2; // @[rvcsr.scala 531:26:@3212.4]
  wire [2:0] _T_1334; // @[rvcsr.scala 514:30:@3193.8]
  wire  dcsr_ebreakh; // @[rvcsr.scala 531:26:@3212.4]
  wire [1:0] _T_1335; // @[rvcsr.scala 514:30:@3194.8]
  wire [3:0] dcsr_xdebugver; // @[rvcsr.scala 531:26:@3212.4]
  wire [11:0] dcsr_rsrvd1; // @[rvcsr.scala 531:26:@3212.4]
  wire [15:0] _T_1336; // @[rvcsr.scala 514:30:@3195.8]
  wire [17:0] _T_1337; // @[rvcsr.scala 514:30:@3196.8]
  wire [20:0] _T_1338; // @[rvcsr.scala 514:30:@3197.8]
  wire [31:0] _T_1339; // @[rvcsr.scala 514:30:@3198.8]
  wire [31:0] _GEN_168; // @[rvcsr.scala 510:38:@3155.6]
  wire [31:0] _GEN_169; // @[rvcsr.scala 517:37:@3201.6]
  wire [31:0] _GEN_170; // @[rvcsr.scala 521:43:@3204.6]
  wire [31:0] _GEN_171; // @[rvcsr.scala 525:43:@3207.6]
  wire [31:0] _GEN_174; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_177; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_178; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_179; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_180; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_181; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_182; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_183; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_186; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_187; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_188; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_189; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_190; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_191; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_192; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_193; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_194; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_195; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_196; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_197; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_198; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_199; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_200; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_201; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_202; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_203; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_204; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_205; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_206; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_207; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_208; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_209; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_210; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_211; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_212; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_213; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_214; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_215; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_216; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_217; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_218; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_219; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_220; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_221; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_222; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_223; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_224; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_225; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_226; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_227; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_228; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_229; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_230; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_231; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_232; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_233; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_234; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_235; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_236; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_237; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_238; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_239; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_240; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_241; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_242; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_243; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_244; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_245; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_246; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_247; // @[rvcsr.scala 393:19:@2545.4]
  wire [63:0] _GEN_248; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_249; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_250; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_253; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_254; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_255; // @[rvcsr.scala 393:19:@2545.4]
  wire [31:0] _GEN_256; // @[rvcsr.scala 393:19:@2545.4]
  wire [1:0] _GEN_257; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_279; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_280; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_281; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_282; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_283; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_284; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_285; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_286; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_287; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_288; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_289; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_290; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_291; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_292; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_293; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_294; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_295; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_296; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_297; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_298; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_299; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_300; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_301; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_302; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_303; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_304; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_305; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_306; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_307; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_308; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_309; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_310; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_311; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_312; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_313; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_314; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_315; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_316; // @[rvcsr.scala 531:26:@3212.4]
  wire [63:0] _GEN_317; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_318; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_319; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_320; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_321; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_322; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_323; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_324; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_325; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_326; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_327; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_328; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_329; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_330; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_331; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_332; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_333; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_334; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_335; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_336; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_337; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_338; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_339; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_340; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_341; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_342; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_343; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_344; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_345; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_346; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_347; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_348; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_349; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_350; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_351; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_366; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_367; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_368; // @[rvcsr.scala 531:26:@3212.4]
  wire [31:0] _GEN_369; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_107 = reg_mcycle[31:0]; // @[rvcsr.scala 253:38:@1594.4]
  assign _T_108 = reg_minstret[63:32]; // @[rvcsr.scala 254:42:@1595.4]
  assign _T_111 = reg_mtime[31:0]; // @[rvcsr.scala 258:36:@1598.4]
  assign _T_112 = reg_mtimecmp[63:32]; // @[rvcsr.scala 259:42:@1599.4]
  assign _T_113 = reg_mtime[63:32]; // @[rvcsr.scala 260:37:@1600.4]
  assign _T_115 = reg_mhpmcounters_0[31:0]; // @[rvcsr.scala 273:73:@1602.4]
  assign _T_116 = reg_mhpmcounters_0[63:32]; // @[rvcsr.scala 274:74:@1603.4]
  assign _T_117 = reg_mhpmcounters_1[31:0]; // @[rvcsr.scala 273:73:@1604.4]
  assign _T_118 = reg_mhpmcounters_1[63:32]; // @[rvcsr.scala 274:74:@1605.4]
  assign _T_119 = reg_mhpmcounters_2[31:0]; // @[rvcsr.scala 273:73:@1606.4]
  assign _T_120 = reg_mhpmcounters_2[63:32]; // @[rvcsr.scala 274:74:@1607.4]
  assign _T_121 = reg_mhpmcounters_3[31:0]; // @[rvcsr.scala 273:73:@1608.4]
  assign _T_122 = reg_mhpmcounters_3[63:32]; // @[rvcsr.scala 274:74:@1609.4]
  assign _T_123 = reg_mhpmcounters_4[31:0]; // @[rvcsr.scala 273:73:@1610.4]
  assign _T_124 = reg_mhpmcounters_4[63:32]; // @[rvcsr.scala 274:74:@1611.4]
  assign _T_125 = reg_mhpmcounters_5[31:0]; // @[rvcsr.scala 273:73:@1612.4]
  assign _T_126 = reg_mhpmcounters_5[63:32]; // @[rvcsr.scala 274:74:@1613.4]
  assign _T_127 = reg_mhpmcounters_6[31:0]; // @[rvcsr.scala 273:73:@1614.4]
  assign _T_128 = reg_mhpmcounters_6[63:32]; // @[rvcsr.scala 274:74:@1615.4]
  assign _T_129 = reg_mhpmcounters_7[31:0]; // @[rvcsr.scala 273:73:@1616.4]
  assign _T_130 = reg_mhpmcounters_7[63:32]; // @[rvcsr.scala 274:74:@1617.4]
  assign _T_131 = reg_mhpmcounters_8[31:0]; // @[rvcsr.scala 273:73:@1618.4]
  assign _T_132 = reg_mhpmcounters_8[63:32]; // @[rvcsr.scala 274:74:@1619.4]
  assign _T_133 = reg_mhpmcounters_9[31:0]; // @[rvcsr.scala 273:73:@1620.4]
  assign _T_134 = reg_mhpmcounters_9[63:32]; // @[rvcsr.scala 274:74:@1621.4]
  assign _T_135 = reg_mhpmcounters_10[31:0]; // @[rvcsr.scala 273:73:@1622.4]
  assign _T_136 = reg_mhpmcounters_10[63:32]; // @[rvcsr.scala 274:74:@1623.4]
  assign _T_137 = reg_mhpmcounters_11[31:0]; // @[rvcsr.scala 273:73:@1624.4]
  assign _T_138 = reg_mhpmcounters_11[63:32]; // @[rvcsr.scala 274:74:@1625.4]
  assign _T_139 = reg_mhpmcounters_12[31:0]; // @[rvcsr.scala 273:73:@1626.4]
  assign _T_140 = reg_mhpmcounters_12[63:32]; // @[rvcsr.scala 274:74:@1627.4]
  assign _T_141 = reg_mhpmcounters_13[31:0]; // @[rvcsr.scala 273:73:@1628.4]
  assign _T_142 = reg_mhpmcounters_13[63:32]; // @[rvcsr.scala 274:74:@1629.4]
  assign _T_143 = reg_mhpmcounters_14[31:0]; // @[rvcsr.scala 273:73:@1630.4]
  assign _T_144 = reg_mhpmcounters_14[63:32]; // @[rvcsr.scala 274:74:@1631.4]
  assign _T_145 = reg_mhpmcounters_15[31:0]; // @[rvcsr.scala 273:73:@1632.4]
  assign _T_146 = reg_mhpmcounters_15[63:32]; // @[rvcsr.scala 274:74:@1633.4]
  assign _T_147 = reg_mhpmcounters_16[31:0]; // @[rvcsr.scala 273:73:@1634.4]
  assign _T_148 = reg_mhpmcounters_16[63:32]; // @[rvcsr.scala 274:74:@1635.4]
  assign _T_149 = reg_mhpmcounters_17[31:0]; // @[rvcsr.scala 273:73:@1636.4]
  assign _T_150 = reg_mhpmcounters_17[63:32]; // @[rvcsr.scala 274:74:@1637.4]
  assign _T_151 = reg_mhpmcounters_18[31:0]; // @[rvcsr.scala 273:73:@1638.4]
  assign _T_152 = reg_mhpmcounters_18[63:32]; // @[rvcsr.scala 274:74:@1639.4]
  assign _T_153 = reg_mhpmcounters_19[31:0]; // @[rvcsr.scala 273:73:@1640.4]
  assign _T_154 = reg_mhpmcounters_19[63:32]; // @[rvcsr.scala 274:74:@1641.4]
  assign _T_155 = reg_mhpmcounters_20[31:0]; // @[rvcsr.scala 273:73:@1642.4]
  assign _T_156 = reg_mhpmcounters_20[63:32]; // @[rvcsr.scala 274:74:@1643.4]
  assign _T_157 = reg_mhpmcounters_21[31:0]; // @[rvcsr.scala 273:73:@1644.4]
  assign _T_158 = reg_mhpmcounters_21[63:32]; // @[rvcsr.scala 274:74:@1645.4]
  assign _T_159 = reg_mhpmcounters_22[31:0]; // @[rvcsr.scala 273:73:@1646.4]
  assign _T_160 = reg_mhpmcounters_22[63:32]; // @[rvcsr.scala 274:74:@1647.4]
  assign _T_161 = reg_mhpmcounters_23[31:0]; // @[rvcsr.scala 273:73:@1648.4]
  assign _T_162 = reg_mhpmcounters_23[63:32]; // @[rvcsr.scala 274:74:@1649.4]
  assign _T_163 = reg_mhpmcounters_24[31:0]; // @[rvcsr.scala 273:73:@1650.4]
  assign _T_164 = reg_mhpmcounters_24[63:32]; // @[rvcsr.scala 274:74:@1651.4]
  assign _T_165 = reg_mhpmcounters_25[31:0]; // @[rvcsr.scala 273:73:@1652.4]
  assign _T_166 = reg_mhpmcounters_25[63:32]; // @[rvcsr.scala 274:74:@1653.4]
  assign _T_167 = reg_mhpmcounters_26[31:0]; // @[rvcsr.scala 273:73:@1654.4]
  assign _T_168 = reg_mhpmcounters_26[63:32]; // @[rvcsr.scala 274:74:@1655.4]
  assign _T_169 = reg_mhpmcounters_27[31:0]; // @[rvcsr.scala 273:73:@1656.4]
  assign _T_170 = reg_mhpmcounters_27[63:32]; // @[rvcsr.scala 274:74:@1657.4]
  assign _T_171 = reg_mhpmcounters_28[31:0]; // @[rvcsr.scala 273:73:@1658.4]
  assign _T_172 = reg_mhpmcounters_28[63:32]; // @[rvcsr.scala 274:74:@1659.4]
  assign counteren_CY = reg_mcounteren[0]; // @[rvcsr.scala 281:48:@1663.4]
  assign counteren_TM = reg_mcounteren[1]; // @[rvcsr.scala 281:48:@1665.4]
  assign counteren_IR = reg_mcounteren[2]; // @[rvcsr.scala 281:48:@1667.4]
  assign counteren_HPM_0 = reg_mcounteren[3]; // @[rvcsr.scala 281:48:@1669.4]
  assign counteren_HPM_1 = reg_mcounteren[4]; // @[rvcsr.scala 281:48:@1671.4]
  assign counteren_HPM_2 = reg_mcounteren[5]; // @[rvcsr.scala 281:48:@1673.4]
  assign counteren_HPM_3 = reg_mcounteren[6]; // @[rvcsr.scala 281:48:@1675.4]
  assign counteren_HPM_4 = reg_mcounteren[7]; // @[rvcsr.scala 281:48:@1677.4]
  assign counteren_HPM_5 = reg_mcounteren[8]; // @[rvcsr.scala 281:48:@1679.4]
  assign counteren_HPM_6 = reg_mcounteren[9]; // @[rvcsr.scala 281:48:@1681.4]
  assign counteren_HPM_7 = reg_mcounteren[10]; // @[rvcsr.scala 281:48:@1683.4]
  assign counteren_HPM_8 = reg_mcounteren[11]; // @[rvcsr.scala 281:48:@1685.4]
  assign counteren_HPM_9 = reg_mcounteren[12]; // @[rvcsr.scala 281:48:@1687.4]
  assign counteren_HPM_10 = reg_mcounteren[13]; // @[rvcsr.scala 281:48:@1689.4]
  assign counteren_HPM_11 = reg_mcounteren[14]; // @[rvcsr.scala 281:48:@1691.4]
  assign counteren_HPM_12 = reg_mcounteren[15]; // @[rvcsr.scala 281:48:@1693.4]
  assign counteren_HPM_13 = reg_mcounteren[16]; // @[rvcsr.scala 281:48:@1695.4]
  assign counteren_HPM_14 = reg_mcounteren[17]; // @[rvcsr.scala 281:48:@1697.4]
  assign counteren_HPM_15 = reg_mcounteren[18]; // @[rvcsr.scala 281:48:@1699.4]
  assign counteren_HPM_16 = reg_mcounteren[19]; // @[rvcsr.scala 281:48:@1701.4]
  assign counteren_HPM_17 = reg_mcounteren[20]; // @[rvcsr.scala 281:48:@1703.4]
  assign counteren_HPM_18 = reg_mcounteren[21]; // @[rvcsr.scala 281:48:@1705.4]
  assign counteren_HPM_19 = reg_mcounteren[22]; // @[rvcsr.scala 281:48:@1707.4]
  assign counteren_HPM_20 = reg_mcounteren[23]; // @[rvcsr.scala 281:48:@1709.4]
  assign counteren_HPM_21 = reg_mcounteren[24]; // @[rvcsr.scala 281:48:@1711.4]
  assign counteren_HPM_22 = reg_mcounteren[25]; // @[rvcsr.scala 281:48:@1713.4]
  assign counteren_HPM_23 = reg_mcounteren[26]; // @[rvcsr.scala 281:48:@1715.4]
  assign counteren_HPM_24 = reg_mcounteren[27]; // @[rvcsr.scala 281:48:@1717.4]
  assign counteren_HPM_25 = reg_mcounteren[28]; // @[rvcsr.scala 281:48:@1719.4]
  assign counteren_HPM_26 = reg_mcounteren[29]; // @[rvcsr.scala 281:48:@1721.4]
  assign counteren_HPM_27 = reg_mcounteren[30]; // @[rvcsr.scala 281:48:@1723.4]
  assign counteren_HPM_28 = reg_mcounteren[31]; // @[rvcsr.scala 281:48:@1725.4]
  assign _T_216 = reg_mcycle + 64'h1; // @[rvcsr.scala 284:34:@1728.6]
  assign _T_217 = _T_216[63:0]; // @[rvcsr.scala 284:34:@1729.6]
  assign _GEN_0 = counteren_CY ? _T_217 : reg_mcycle; // @[rvcsr.scala 283:24:@1727.4]
  assign _T_219 = reg_mtime + 64'h1; // @[rvcsr.scala 288:32:@1733.6]
  assign _T_220 = _T_219[63:0]; // @[rvcsr.scala 288:32:@1734.6]
  assign _GEN_1 = counteren_TM ? _T_220 : reg_mtime; // @[rvcsr.scala 287:24:@1732.4]
  assign _T_222 = reg_minstret + 64'h1; // @[rvcsr.scala 292:38:@1738.6]
  assign _T_223 = _T_222[63:0]; // @[rvcsr.scala 292:38:@1739.6]
  assign _GEN_2 = counteren_IR ? _T_223 : reg_minstret; // @[rvcsr.scala 291:24:@1737.4]
  assign _T_225 = reg_mhpmcounters_0 + 64'h1; // @[rvcsr.scala 297:56:@1743.6]
  assign _T_226 = _T_225[63:0]; // @[rvcsr.scala 297:56:@1744.6]
  assign _GEN_3 = counteren_HPM_0 ? _T_226 : reg_mhpmcounters_0; // @[rvcsr.scala 296:32:@1742.4]
  assign _T_228 = reg_mhpmcounters_1 + 64'h1; // @[rvcsr.scala 297:56:@1748.6]
  assign _T_229 = _T_228[63:0]; // @[rvcsr.scala 297:56:@1749.6]
  assign _GEN_4 = counteren_HPM_1 ? _T_229 : reg_mhpmcounters_1; // @[rvcsr.scala 296:32:@1747.4]
  assign _T_231 = reg_mhpmcounters_2 + 64'h1; // @[rvcsr.scala 297:56:@1753.6]
  assign _T_232 = _T_231[63:0]; // @[rvcsr.scala 297:56:@1754.6]
  assign _GEN_5 = counteren_HPM_2 ? _T_232 : reg_mhpmcounters_2; // @[rvcsr.scala 296:32:@1752.4]
  assign _T_234 = reg_mhpmcounters_3 + 64'h1; // @[rvcsr.scala 297:56:@1758.6]
  assign _T_235 = _T_234[63:0]; // @[rvcsr.scala 297:56:@1759.6]
  assign _GEN_6 = counteren_HPM_3 ? _T_235 : reg_mhpmcounters_3; // @[rvcsr.scala 296:32:@1757.4]
  assign _T_237 = reg_mhpmcounters_4 + 64'h1; // @[rvcsr.scala 297:56:@1763.6]
  assign _T_238 = _T_237[63:0]; // @[rvcsr.scala 297:56:@1764.6]
  assign _GEN_7 = counteren_HPM_4 ? _T_238 : reg_mhpmcounters_4; // @[rvcsr.scala 296:32:@1762.4]
  assign _T_240 = reg_mhpmcounters_5 + 64'h1; // @[rvcsr.scala 297:56:@1768.6]
  assign _T_241 = _T_240[63:0]; // @[rvcsr.scala 297:56:@1769.6]
  assign _GEN_8 = counteren_HPM_5 ? _T_241 : reg_mhpmcounters_5; // @[rvcsr.scala 296:32:@1767.4]
  assign _T_243 = reg_mhpmcounters_6 + 64'h1; // @[rvcsr.scala 297:56:@1773.6]
  assign _T_244 = _T_243[63:0]; // @[rvcsr.scala 297:56:@1774.6]
  assign _GEN_9 = counteren_HPM_6 ? _T_244 : reg_mhpmcounters_6; // @[rvcsr.scala 296:32:@1772.4]
  assign _T_246 = reg_mhpmcounters_7 + 64'h1; // @[rvcsr.scala 297:56:@1778.6]
  assign _T_247 = _T_246[63:0]; // @[rvcsr.scala 297:56:@1779.6]
  assign _GEN_10 = counteren_HPM_7 ? _T_247 : reg_mhpmcounters_7; // @[rvcsr.scala 296:32:@1777.4]
  assign _T_249 = reg_mhpmcounters_8 + 64'h1; // @[rvcsr.scala 297:56:@1783.6]
  assign _T_250 = _T_249[63:0]; // @[rvcsr.scala 297:56:@1784.6]
  assign _GEN_11 = counteren_HPM_8 ? _T_250 : reg_mhpmcounters_8; // @[rvcsr.scala 296:32:@1782.4]
  assign _T_252 = reg_mhpmcounters_9 + 64'h1; // @[rvcsr.scala 297:56:@1788.6]
  assign _T_253 = _T_252[63:0]; // @[rvcsr.scala 297:56:@1789.6]
  assign _GEN_12 = counteren_HPM_9 ? _T_253 : reg_mhpmcounters_9; // @[rvcsr.scala 296:32:@1787.4]
  assign _T_255 = reg_mhpmcounters_10 + 64'h1; // @[rvcsr.scala 297:56:@1793.6]
  assign _T_256 = _T_255[63:0]; // @[rvcsr.scala 297:56:@1794.6]
  assign _GEN_13 = counteren_HPM_10 ? _T_256 : reg_mhpmcounters_10; // @[rvcsr.scala 296:32:@1792.4]
  assign _T_258 = reg_mhpmcounters_11 + 64'h1; // @[rvcsr.scala 297:56:@1798.6]
  assign _T_259 = _T_258[63:0]; // @[rvcsr.scala 297:56:@1799.6]
  assign _GEN_14 = counteren_HPM_11 ? _T_259 : reg_mhpmcounters_11; // @[rvcsr.scala 296:32:@1797.4]
  assign _T_261 = reg_mhpmcounters_12 + 64'h1; // @[rvcsr.scala 297:56:@1803.6]
  assign _T_262 = _T_261[63:0]; // @[rvcsr.scala 297:56:@1804.6]
  assign _GEN_15 = counteren_HPM_12 ? _T_262 : reg_mhpmcounters_12; // @[rvcsr.scala 296:32:@1802.4]
  assign _T_264 = reg_mhpmcounters_13 + 64'h1; // @[rvcsr.scala 297:56:@1808.6]
  assign _T_265 = _T_264[63:0]; // @[rvcsr.scala 297:56:@1809.6]
  assign _GEN_16 = counteren_HPM_13 ? _T_265 : reg_mhpmcounters_13; // @[rvcsr.scala 296:32:@1807.4]
  assign _T_267 = reg_mhpmcounters_14 + 64'h1; // @[rvcsr.scala 297:56:@1813.6]
  assign _T_268 = _T_267[63:0]; // @[rvcsr.scala 297:56:@1814.6]
  assign _GEN_17 = counteren_HPM_14 ? _T_268 : reg_mhpmcounters_14; // @[rvcsr.scala 296:32:@1812.4]
  assign _T_270 = reg_mhpmcounters_15 + 64'h1; // @[rvcsr.scala 297:56:@1818.6]
  assign _T_271 = _T_270[63:0]; // @[rvcsr.scala 297:56:@1819.6]
  assign _GEN_18 = counteren_HPM_15 ? _T_271 : reg_mhpmcounters_15; // @[rvcsr.scala 296:32:@1817.4]
  assign _T_273 = reg_mhpmcounters_16 + 64'h1; // @[rvcsr.scala 297:56:@1823.6]
  assign _T_274 = _T_273[63:0]; // @[rvcsr.scala 297:56:@1824.6]
  assign _GEN_19 = counteren_HPM_16 ? _T_274 : reg_mhpmcounters_16; // @[rvcsr.scala 296:32:@1822.4]
  assign _T_276 = reg_mhpmcounters_17 + 64'h1; // @[rvcsr.scala 297:56:@1828.6]
  assign _T_277 = _T_276[63:0]; // @[rvcsr.scala 297:56:@1829.6]
  assign _GEN_20 = counteren_HPM_17 ? _T_277 : reg_mhpmcounters_17; // @[rvcsr.scala 296:32:@1827.4]
  assign _T_279 = reg_mhpmcounters_18 + 64'h1; // @[rvcsr.scala 297:56:@1833.6]
  assign _T_280 = _T_279[63:0]; // @[rvcsr.scala 297:56:@1834.6]
  assign _GEN_21 = counteren_HPM_18 ? _T_280 : reg_mhpmcounters_18; // @[rvcsr.scala 296:32:@1832.4]
  assign _T_282 = reg_mhpmcounters_19 + 64'h1; // @[rvcsr.scala 297:56:@1838.6]
  assign _T_283 = _T_282[63:0]; // @[rvcsr.scala 297:56:@1839.6]
  assign _GEN_22 = counteren_HPM_19 ? _T_283 : reg_mhpmcounters_19; // @[rvcsr.scala 296:32:@1837.4]
  assign _T_285 = reg_mhpmcounters_20 + 64'h1; // @[rvcsr.scala 297:56:@1843.6]
  assign _T_286 = _T_285[63:0]; // @[rvcsr.scala 297:56:@1844.6]
  assign _GEN_23 = counteren_HPM_20 ? _T_286 : reg_mhpmcounters_20; // @[rvcsr.scala 296:32:@1842.4]
  assign _T_288 = reg_mhpmcounters_21 + 64'h1; // @[rvcsr.scala 297:56:@1848.6]
  assign _T_289 = _T_288[63:0]; // @[rvcsr.scala 297:56:@1849.6]
  assign _GEN_24 = counteren_HPM_21 ? _T_289 : reg_mhpmcounters_21; // @[rvcsr.scala 296:32:@1847.4]
  assign _T_291 = reg_mhpmcounters_22 + 64'h1; // @[rvcsr.scala 297:56:@1853.6]
  assign _T_292 = _T_291[63:0]; // @[rvcsr.scala 297:56:@1854.6]
  assign _GEN_25 = counteren_HPM_22 ? _T_292 : reg_mhpmcounters_22; // @[rvcsr.scala 296:32:@1852.4]
  assign _T_294 = reg_mhpmcounters_23 + 64'h1; // @[rvcsr.scala 297:56:@1858.6]
  assign _T_295 = _T_294[63:0]; // @[rvcsr.scala 297:56:@1859.6]
  assign _GEN_26 = counteren_HPM_23 ? _T_295 : reg_mhpmcounters_23; // @[rvcsr.scala 296:32:@1857.4]
  assign _T_297 = reg_mhpmcounters_24 + 64'h1; // @[rvcsr.scala 297:56:@1863.6]
  assign _T_298 = _T_297[63:0]; // @[rvcsr.scala 297:56:@1864.6]
  assign _GEN_27 = counteren_HPM_24 ? _T_298 : reg_mhpmcounters_24; // @[rvcsr.scala 296:32:@1862.4]
  assign _T_300 = reg_mhpmcounters_25 + 64'h1; // @[rvcsr.scala 297:56:@1868.6]
  assign _T_301 = _T_300[63:0]; // @[rvcsr.scala 297:56:@1869.6]
  assign _GEN_28 = counteren_HPM_25 ? _T_301 : reg_mhpmcounters_25; // @[rvcsr.scala 296:32:@1867.4]
  assign _T_303 = reg_mhpmcounters_26 + 64'h1; // @[rvcsr.scala 297:56:@1873.6]
  assign _T_304 = _T_303[63:0]; // @[rvcsr.scala 297:56:@1874.6]
  assign _GEN_29 = counteren_HPM_26 ? _T_304 : reg_mhpmcounters_26; // @[rvcsr.scala 296:32:@1872.4]
  assign _T_306 = reg_mhpmcounters_27 + 64'h1; // @[rvcsr.scala 297:56:@1878.6]
  assign _T_307 = _T_306[63:0]; // @[rvcsr.scala 297:56:@1879.6]
  assign _GEN_30 = counteren_HPM_27 ? _T_307 : reg_mhpmcounters_27; // @[rvcsr.scala 296:32:@1877.4]
  assign _T_309 = reg_mhpmcounters_28 + 64'h1; // @[rvcsr.scala 297:56:@1883.6]
  assign _T_310 = _T_309[63:0]; // @[rvcsr.scala 297:56:@1884.6]
  assign _GEN_31 = counteren_HPM_28 ? _T_310 : reg_mhpmcounters_28; // @[rvcsr.scala 296:32:@1882.4]
  assign _T_318 = reg_mstatus[0]; // @[rvcsr.scala 311:40:@1893.4]
  assign _T_319 = reg_mstatus[1]; // @[rvcsr.scala 311:40:@1895.4]
  assign _T_320 = reg_mstatus[2]; // @[rvcsr.scala 311:40:@1897.4]
  assign _T_321 = reg_mstatus[3]; // @[rvcsr.scala 311:40:@1899.4]
  assign _T_322 = reg_mstatus[4]; // @[rvcsr.scala 311:40:@1901.4]
  assign _T_323 = reg_mstatus[5]; // @[rvcsr.scala 311:40:@1903.4]
  assign _T_324 = reg_mstatus[6]; // @[rvcsr.scala 311:40:@1905.4]
  assign _T_325 = reg_mstatus[7]; // @[rvcsr.scala 311:40:@1907.4]
  assign _T_326 = reg_mstatus[8]; // @[rvcsr.scala 311:40:@1909.4]
  assign _T_327 = reg_mstatus[10:9]; // @[rvcsr.scala 311:40:@1911.4]
  assign _T_328 = reg_mstatus[12:11]; // @[rvcsr.scala 311:40:@1913.4]
  assign _T_329 = reg_mstatus[14:13]; // @[rvcsr.scala 311:40:@1915.4]
  assign _T_330 = reg_mstatus[16:15]; // @[rvcsr.scala 311:40:@1917.4]
  assign _T_331 = reg_mstatus[17]; // @[rvcsr.scala 311:40:@1919.4]
  assign _T_332 = reg_mstatus[18]; // @[rvcsr.scala 311:40:@1921.4]
  assign _T_333 = reg_mstatus[19]; // @[rvcsr.scala 311:40:@1923.4]
  assign _T_334 = reg_mstatus[20]; // @[rvcsr.scala 311:40:@1925.4]
  assign _T_335 = reg_mstatus[21]; // @[rvcsr.scala 311:40:@1927.4]
  assign _T_336 = reg_mstatus[22]; // @[rvcsr.scala 311:40:@1929.4]
  assign _T_337 = reg_mstatus[30:23]; // @[rvcsr.scala 311:40:@1931.4]
  assign _T_338 = reg_mstatus[31]; // @[rvcsr.scala 311:40:@1933.4]
  assign _T_344 = reg_mie[30:0]; // @[:@1958.4]
  assign mie_USIE = _T_344[0]; // @[rvcsr.scala 313:32:@1960.4]
  assign mie_SSIE = _T_344[1]; // @[rvcsr.scala 313:32:@1962.4]
  assign mie_rsrvd4 = _T_344[2]; // @[rvcsr.scala 313:32:@1964.4]
  assign _T_348 = _T_344[3]; // @[rvcsr.scala 313:32:@1966.4]
  assign mie_UTIE = _T_344[4]; // @[rvcsr.scala 313:32:@1968.4]
  assign mie_STIE = _T_344[5]; // @[rvcsr.scala 313:32:@1970.4]
  assign mie_rsrvd3 = _T_344[6]; // @[rvcsr.scala 313:32:@1972.4]
  assign _T_352 = _T_344[7]; // @[rvcsr.scala 313:32:@1974.4]
  assign mie_UEIE = _T_344[8]; // @[rvcsr.scala 313:32:@1976.4]
  assign mie_SEIE = _T_344[9]; // @[rvcsr.scala 313:32:@1978.4]
  assign mie_rsrvd2 = _T_344[10]; // @[rvcsr.scala 313:32:@1980.4]
  assign mie_MEIE = _T_344[11]; // @[rvcsr.scala 313:32:@1982.4]
  assign mie_rsrvd1 = _T_344[30:12]; // @[rvcsr.scala 313:32:@1984.4]
  assign _T_363 = reg_mip[30:0]; // @[:@2001.4]
  assign mip_USIP = _T_363[0]; // @[rvcsr.scala 315:32:@2003.4]
  assign mip_SSIP = _T_363[1]; // @[rvcsr.scala 315:32:@2005.4]
  assign mip_rsrvd4 = _T_363[2]; // @[rvcsr.scala 315:32:@2007.4]
  assign _T_367 = _T_363[3]; // @[rvcsr.scala 315:32:@2009.4]
  assign mip_UTIP = _T_363[4]; // @[rvcsr.scala 315:32:@2011.4]
  assign mip_STIP = _T_363[5]; // @[rvcsr.scala 315:32:@2013.4]
  assign mip_rsrvd3 = _T_363[6]; // @[rvcsr.scala 315:32:@2015.4]
  assign _T_371 = _T_363[7]; // @[rvcsr.scala 315:32:@2017.4]
  assign mip_UEIP = _T_363[8]; // @[rvcsr.scala 315:32:@2019.4]
  assign mip_SEIP = _T_363[9]; // @[rvcsr.scala 315:32:@2021.4]
  assign mip_rsrvd2 = _T_363[10]; // @[rvcsr.scala 315:32:@2023.4]
  assign mip_MEIP = _T_363[11]; // @[rvcsr.scala 315:32:@2025.4]
  assign mip_rsrvd1 = _T_363[30:12]; // @[rvcsr.scala 315:32:@2027.4]
  assign _T_383 = reg_dcsr[1:0]; // @[rvcsr.scala 317:34:@2046.4]
  assign _T_384 = reg_dcsr[2]; // @[rvcsr.scala 317:34:@2048.4]
  assign _T_385 = reg_dcsr[5:3]; // @[rvcsr.scala 317:34:@2050.4]
  assign _T_386 = reg_dcsr[8:6]; // @[rvcsr.scala 317:34:@2052.4]
  assign _T_387 = reg_dcsr[9]; // @[rvcsr.scala 317:34:@2054.4]
  assign _T_388 = reg_dcsr[10]; // @[rvcsr.scala 317:34:@2056.4]
  assign _T_389 = reg_dcsr[11]; // @[rvcsr.scala 317:34:@2058.4]
  assign _T_390 = reg_dcsr[12]; // @[rvcsr.scala 317:34:@2060.4]
  assign _T_391 = reg_dcsr[13]; // @[rvcsr.scala 317:34:@2062.4]
  assign _T_392 = reg_dcsr[14]; // @[rvcsr.scala 317:34:@2064.4]
  assign _T_393 = reg_dcsr[15]; // @[rvcsr.scala 317:34:@2066.4]
  assign _T_394 = reg_dcsr[27:16]; // @[rvcsr.scala 317:34:@2068.4]
  assign _T_395 = reg_dcsr[31:28]; // @[rvcsr.scala 317:34:@2070.4]
  assign csr_priv = io_addr[9:8]; // @[rvcsr.scala 319:27:@2085.4]
  assign legal_priv = reg_priv >= csr_priv; // @[rvcsr.scala 320:28:@2086.4]
  assign priv_inst = io_op == 3'h4; // @[rvcsr.scala 321:28:@2087.4]
  assign priv_inst_type = io_addr[2:0]; // @[rvcsr.scala 322:33:@2088.4]
  assign _T_396 = legal_priv & priv_inst; // @[rvcsr.scala 323:33:@2089.4]
  assign _T_398 = priv_inst_type == 3'h0; // @[rvcsr.scala 323:61:@2090.4]
  assign inst_ecall = _T_396 & _T_398; // @[rvcsr.scala 323:44:@2091.4]
  assign _T_401 = priv_inst_type == 3'h1; // @[rvcsr.scala 324:62:@2093.4]
  assign inst_ebreak = _T_396 & _T_401; // @[rvcsr.scala 324:45:@2094.4]
  assign _T_404 = priv_inst_type == 3'h2; // @[rvcsr.scala 325:59:@2096.4]
  assign inst_ret = _T_396 & _T_404; // @[rvcsr.scala 325:42:@2097.4]
  assign _T_405 = inst_ecall | inst_ebreak; // @[rvcsr.scala 328:31:@2098.4]
  assign _T_406 = _T_405 | inst_ret; // @[rvcsr.scala 328:45:@2099.4]
  assign _T_407 = reg_mtime >= reg_mtimecmp; // @[rvcsr.scala 331:21:@2101.4]
  assign _T_409 = {mip_rsrvd4,mip_SSIP}; // @[rvcsr.scala 333:24:@2104.6]
  assign _T_410 = {_T_409,mip_USIP}; // @[rvcsr.scala 333:24:@2105.6]
  assign _T_411 = {mip_STIP,mip_UTIP}; // @[rvcsr.scala 333:24:@2106.6]
  assign _T_690 = io_addr[11]; // @[rvcsr.scala 382:28:@2294.4]
  assign _T_691 = io_addr[10]; // @[rvcsr.scala 382:40:@2295.4]
  assign read_only = _T_690 & _T_691; // @[rvcsr.scala 382:32:@2296.4]
  assign _T_693 = read_only == 1'h0; // @[rvcsr.scala 384:20:@2298.4]
  assign _T_695 = priv_inst == 1'h0; // @[rvcsr.scala 384:33:@2299.4]
  assign _T_696 = _T_693 & _T_695; // @[rvcsr.scala 384:31:@2300.4]
  assign csr_wen = _T_696 & legal_priv; // @[rvcsr.scala 384:43:@2301.4]
  assign _T_491 = io_addr == 12'h344; // @[rvcsr.scala 380:61:@2194.4]
  assign _T_1046 = io_op != 3'h1; // @[rvcsr.scala 392:30:@2535.4]
  assign _T_1048 = _T_1046 ? io_rdata : 32'h0; // @[rvcsr.scala 392:22:@2536.4]
  assign _T_1049 = io_op != 3'h3; // @[rvcsr.scala 392:73:@2537.4]
  assign _T_1051 = _T_1049 ? io_wdata : 32'h0; // @[rvcsr.scala 392:65:@2538.4]
  assign _T_1052 = _T_1048 | _T_1051; // @[rvcsr.scala 392:60:@2539.4]
  assign _T_1053 = io_op == 3'h3; // @[rvcsr.scala 392:119:@2540.4]
  assign _T_1055 = _T_1053 ? io_wdata : 32'h0; // @[rvcsr.scala 392:111:@2541.4]
  assign _T_1056 = ~ _T_1055; // @[rvcsr.scala 392:107:@2542.4]
  assign csr_wdata = _T_1052 & _T_1056; // @[rvcsr.scala 392:104:@2543.4]
  assign _T_1152 = csr_wdata[30:0]; // @[:@2688.8]
  assign _T_1156 = _T_1152[3]; // @[rvcsr.scala 435:47:@2696.8]
  assign _GEN_67 = _T_491 ? _T_1156 : _T_367; // @[rvcsr.scala 434:37:@2686.6]
  assign mip_MSIP = csr_wen ? _GEN_67 : _T_367; // @[rvcsr.scala 393:19:@2545.4]
  assign _T_412 = {_T_411,mip_MSIP}; // @[rvcsr.scala 333:24:@2107.6]
  assign _T_413 = {_T_412,_T_410}; // @[rvcsr.scala 333:24:@2108.6]
  assign _T_1160 = _T_1152[7]; // @[rvcsr.scala 435:47:@2704.8]
  assign _GEN_32 = _T_407 ? 1'h1 : _T_371; // @[rvcsr.scala 331:38:@2102.4]
  assign _GEN_66 = _T_491 ? _T_1160 : _GEN_32; // @[rvcsr.scala 434:37:@2686.6]
  assign mip_MTIP = csr_wen ? _GEN_66 : _GEN_32; // @[rvcsr.scala 393:19:@2545.4]
  assign _T_414 = {mip_UEIP,mip_MTIP}; // @[rvcsr.scala 333:24:@2109.6]
  assign _T_415 = {_T_414,mip_rsrvd3}; // @[rvcsr.scala 333:24:@2110.6]
  assign _T_416 = {mip_rsrvd2,mip_SEIP}; // @[rvcsr.scala 333:24:@2111.6]
  assign _T_417 = {mip_rsrvd1,mip_MEIP}; // @[rvcsr.scala 333:24:@2112.6]
  assign _T_418 = {_T_417,_T_416}; // @[rvcsr.scala 333:24:@2113.6]
  assign _T_419 = {_T_418,_T_415}; // @[rvcsr.scala 333:24:@2114.6]
  assign _T_420 = {_T_419,_T_413}; // @[rvcsr.scala 333:24:@2115.6]
  assign _GEN_33 = _T_407 ? {{1'd0}, _T_420} : reg_mip; // @[rvcsr.scala 331:38:@2102.4]
  assign _T_421 = csr_priv == 2'h3; // @[rvcsr.scala 337:32:@2118.4]
  assign _T_422 = inst_ret & _T_421; // @[rvcsr.scala 337:20:@2119.4]
  assign _T_425 = _T_691 == 1'h0; // @[rvcsr.scala 337:61:@2121.4]
  assign _T_426 = _T_422 & _T_425; // @[rvcsr.scala 337:46:@2122.4]
  assign mstatus_SIE = reset ? 1'h0 : _T_319; // @[rvcsr.scala 531:26:@3212.4]
  assign mstatus_UIE = reset ? 1'h0 : _T_318; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_428 = {mstatus_SIE,mstatus_UIE}; // @[rvcsr.scala 342:32:@2128.6]
  assign mstatus_UPIE = reset ? 1'h0 : _T_322; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_469 = io_addr == 12'h300; // @[rvcsr.scala 380:61:@2183.4]
  assign _T_1066 = csr_wdata[3]; // @[rvcsr.scala 396:55:@2556.8]
  assign _T_1070 = csr_wdata[7]; // @[rvcsr.scala 396:55:@2564.8]
  assign _GEN_35 = _T_426 ? 1'h1 : _T_325; // @[rvcsr.scala 337:73:@2123.4]
  assign _GEN_55 = _T_469 ? _T_1070 : _GEN_35; // @[rvcsr.scala 395:41:@2546.6]
  assign _GEN_173 = csr_wen ? _GEN_55 : _GEN_35; // @[rvcsr.scala 393:19:@2545.4]
  assign mstatus_MPIE = reset ? 1'h0 : _GEN_173; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_34 = _T_426 ? mstatus_MPIE : _T_321; // @[rvcsr.scala 337:73:@2123.4]
  assign _GEN_54 = _T_469 ? _T_1066 : _GEN_34; // @[rvcsr.scala 395:41:@2546.6]
  assign _GEN_172 = csr_wen ? _GEN_54 : _GEN_34; // @[rvcsr.scala 393:19:@2545.4]
  assign mstatus_MIE = reset ? 1'h0 : _GEN_172; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_429 = {mstatus_UPIE,mstatus_MIE}; // @[rvcsr.scala 342:32:@2129.6]
  assign mstatus_rsrvd4 = reset ? 1'h0 : _T_320; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_430 = {_T_429,mstatus_rsrvd4}; // @[rvcsr.scala 342:32:@2130.6]
  assign _T_431 = {_T_430,_T_428}; // @[rvcsr.scala 342:32:@2131.6]
  assign mstatus_rsrvd3 = reset ? 1'h0 : _T_324; // @[rvcsr.scala 531:26:@3212.4]
  assign mstatus_SPIE = reset ? 1'h0 : _T_323; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_432 = {mstatus_rsrvd3,mstatus_SPIE}; // @[rvcsr.scala 342:32:@2132.6]
  assign mstatus_rsrvd2 = reset ? 2'h0 : _T_327; // @[rvcsr.scala 531:26:@3212.4]
  assign mstatus_SPP = reset ? 1'h0 : _T_326; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_433 = {mstatus_rsrvd2,mstatus_SPP}; // @[rvcsr.scala 342:32:@2133.6]
  assign _T_434 = {_T_433,mstatus_MPIE}; // @[rvcsr.scala 342:32:@2134.6]
  assign _T_435 = {_T_434,_T_432}; // @[rvcsr.scala 342:32:@2135.6]
  assign _T_436 = {_T_435,_T_431}; // @[rvcsr.scala 342:32:@2136.6]
  assign mstatus_FS = reset ? 2'h0 : _T_329; // @[rvcsr.scala 531:26:@3212.4]
  assign mstatus_MPP = reset ? 2'h3 : _T_328; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_437 = {mstatus_FS,mstatus_MPP}; // @[rvcsr.scala 342:32:@2137.6]
  assign mstatus_SUM = reset ? 1'h0 : _T_332; // @[rvcsr.scala 531:26:@3212.4]
  assign mstatus_MPRV = reset ? 1'h0 : _T_331; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_438 = {mstatus_SUM,mstatus_MPRV}; // @[rvcsr.scala 342:32:@2138.6]
  assign mstatus_XS = reset ? 2'h0 : _T_330; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_439 = {_T_438,mstatus_XS}; // @[rvcsr.scala 342:32:@2139.6]
  assign _T_440 = {_T_439,_T_437}; // @[rvcsr.scala 342:32:@2140.6]
  assign mstatus_TW = reset ? 1'h0 : _T_335; // @[rvcsr.scala 531:26:@3212.4]
  assign mstatus_TVM = reset ? 1'h0 : _T_334; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_441 = {mstatus_TW,mstatus_TVM}; // @[rvcsr.scala 342:32:@2141.6]
  assign mstatus_MXR = reset ? 1'h0 : _T_333; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_442 = {_T_441,mstatus_MXR}; // @[rvcsr.scala 342:32:@2142.6]
  assign mstatus_SD = reset ? 1'h0 : _T_338; // @[rvcsr.scala 531:26:@3212.4]
  assign mstatus_rsrvd1 = reset ? 8'h0 : _T_337; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_443 = {mstatus_SD,mstatus_rsrvd1}; // @[rvcsr.scala 342:32:@2143.6]
  assign mstatus_TSR = reset ? 1'h0 : _T_336; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_444 = {_T_443,mstatus_TSR}; // @[rvcsr.scala 342:32:@2144.6]
  assign _T_445 = {_T_444,_T_442}; // @[rvcsr.scala 342:32:@2145.6]
  assign _T_446 = {_T_445,_T_440}; // @[rvcsr.scala 342:32:@2146.6]
  assign _T_447 = {_T_446,_T_436}; // @[rvcsr.scala 342:32:@2147.6]
  assign _GEN_36 = _T_426 ? mstatus_MPP : reg_priv; // @[rvcsr.scala 337:73:@2123.4]
  assign _GEN_38 = _T_426 ? _T_447 : reg_mstatus; // @[rvcsr.scala 337:73:@2123.4]
  assign _GEN_39 = inst_ecall ? 32'hb : reg_mcause; // @[rvcsr.scala 346:21:@2150.4]
  assign _GEN_40 = inst_ecall ? 32'h80000004 : reg_mepc; // @[rvcsr.scala 346:21:@2150.4]
  assign _T_509 = io_addr == 12'h7b0; // @[rvcsr.scala 380:61:@2203.4]
  assign _T_1325 = csr_wdata[15]; // @[rvcsr.scala 511:49:@3179.8]
  assign _GEN_167 = _T_509 ? _T_1325 : _T_393; // @[rvcsr.scala 510:38:@3155.6]
  assign _GEN_252 = csr_wen ? _GEN_167 : _T_393; // @[rvcsr.scala 393:19:@2545.4]
  assign dcsr_ebreakm = reset ? 1'h0 : _GEN_252; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_42 = inst_ebreak ? 32'h3 : _GEN_39; // @[rvcsr.scala 352:22:@2154.4]
  assign _GEN_43 = inst_ebreak ? 32'h80000004 : _GEN_40; // @[rvcsr.scala 352:22:@2154.4]
  assign _T_456 = _T_422 & _T_691; // @[rvcsr.scala 361:46:@2165.4]
  assign dcsr_prv = reset ? 2'h3 : _T_383; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_46 = _T_456 ? dcsr_prv : _GEN_36; // @[rvcsr.scala 361:72:@2166.4]
  assign _GEN_47 = _T_456 ? reg_dpc : _GEN_43; // @[rvcsr.scala 361:72:@2166.4]
  assign _T_458 = 4'h2 == io_core_cause; // @[Conditional.scala 37:30:@2172.6]
  assign _GEN_48 = _T_458 ? {{28'd0}, io_core_cause} : _GEN_42; // @[Conditional.scala 40:58:@2173.6]
  assign _GEN_49 = _T_458 ? io_core_pc : reg_mepc; // @[Conditional.scala 40:58:@2173.6]
  assign _GEN_50 = _T_458 ? 32'h80000004 : _GEN_47; // @[Conditional.scala 40:58:@2173.6]
  assign _GEN_51 = io_core_excp ? _GEN_48 : _GEN_42; // @[rvcsr.scala 368:25:@2171.4]
  assign _GEN_52 = io_core_excp ? _GEN_49 : reg_mepc; // @[rvcsr.scala 368:25:@2171.4]
  assign _GEN_53 = io_core_excp ? _GEN_50 : _GEN_47; // @[rvcsr.scala 368:25:@2171.4]
  assign _T_473 = io_addr == 12'h302; // @[rvcsr.scala 380:61:@2185.4]
  assign _T_475 = io_addr == 12'h303; // @[rvcsr.scala 380:61:@2186.4]
  assign _T_477 = io_addr == 12'h304; // @[rvcsr.scala 380:61:@2187.4]
  assign _T_479 = io_addr == 12'h305; // @[rvcsr.scala 380:61:@2188.4]
  assign _T_481 = io_addr == 12'h306; // @[rvcsr.scala 380:61:@2189.4]
  assign _T_483 = io_addr == 12'h340; // @[rvcsr.scala 380:61:@2190.4]
  assign _T_485 = io_addr == 12'h341; // @[rvcsr.scala 380:61:@2191.4]
  assign _T_487 = io_addr == 12'h342; // @[rvcsr.scala 380:61:@2192.4]
  assign _T_489 = io_addr == 12'h343; // @[rvcsr.scala 380:61:@2193.4]
  assign _T_493 = io_addr == 12'hb00; // @[rvcsr.scala 380:61:@2195.4]
  assign _T_495 = io_addr == 12'hb02; // @[rvcsr.scala 380:61:@2196.4]
  assign _T_497 = io_addr == 12'hb80; // @[rvcsr.scala 380:61:@2197.4]
  assign _T_499 = io_addr == 12'hb82; // @[rvcsr.scala 380:61:@2198.4]
  assign _T_501 = io_addr == 12'hb01; // @[rvcsr.scala 380:61:@2199.4]
  assign _T_503 = io_addr == 12'hb20; // @[rvcsr.scala 380:61:@2200.4]
  assign _T_505 = io_addr == 12'hb81; // @[rvcsr.scala 380:61:@2201.4]
  assign _T_507 = io_addr == 12'hba0; // @[rvcsr.scala 380:61:@2202.4]
  assign _T_511 = io_addr == 12'h7b1; // @[rvcsr.scala 380:61:@2204.4]
  assign _T_513 = io_addr == 12'h7b2; // @[rvcsr.scala 380:61:@2205.4]
  assign _T_515 = io_addr == 12'h7b3; // @[rvcsr.scala 380:61:@2206.4]
  assign _T_517 = io_addr == 12'hb03; // @[rvcsr.scala 380:61:@2207.4]
  assign _T_519 = io_addr == 12'hb83; // @[rvcsr.scala 380:61:@2208.4]
  assign _T_521 = io_addr == 12'hb04; // @[rvcsr.scala 380:61:@2209.4]
  assign _T_523 = io_addr == 12'hb84; // @[rvcsr.scala 380:61:@2210.4]
  assign _T_525 = io_addr == 12'hb05; // @[rvcsr.scala 380:61:@2211.4]
  assign _T_527 = io_addr == 12'hb85; // @[rvcsr.scala 380:61:@2212.4]
  assign _T_529 = io_addr == 12'hb06; // @[rvcsr.scala 380:61:@2213.4]
  assign _T_531 = io_addr == 12'hb86; // @[rvcsr.scala 380:61:@2214.4]
  assign _T_533 = io_addr == 12'hb07; // @[rvcsr.scala 380:61:@2215.4]
  assign _T_535 = io_addr == 12'hb87; // @[rvcsr.scala 380:61:@2216.4]
  assign _T_537 = io_addr == 12'hb08; // @[rvcsr.scala 380:61:@2217.4]
  assign _T_539 = io_addr == 12'hb88; // @[rvcsr.scala 380:61:@2218.4]
  assign _T_541 = io_addr == 12'hb09; // @[rvcsr.scala 380:61:@2219.4]
  assign _T_543 = io_addr == 12'hb89; // @[rvcsr.scala 380:61:@2220.4]
  assign _T_545 = io_addr == 12'hb0a; // @[rvcsr.scala 380:61:@2221.4]
  assign _T_547 = io_addr == 12'hb8a; // @[rvcsr.scala 380:61:@2222.4]
  assign _T_549 = io_addr == 12'hb0b; // @[rvcsr.scala 380:61:@2223.4]
  assign _T_551 = io_addr == 12'hb8b; // @[rvcsr.scala 380:61:@2224.4]
  assign _T_553 = io_addr == 12'hb0c; // @[rvcsr.scala 380:61:@2225.4]
  assign _T_555 = io_addr == 12'hb8c; // @[rvcsr.scala 380:61:@2226.4]
  assign _T_557 = io_addr == 12'hb0d; // @[rvcsr.scala 380:61:@2227.4]
  assign _T_559 = io_addr == 12'hb8d; // @[rvcsr.scala 380:61:@2228.4]
  assign _T_561 = io_addr == 12'hb0e; // @[rvcsr.scala 380:61:@2229.4]
  assign _T_563 = io_addr == 12'hb8e; // @[rvcsr.scala 380:61:@2230.4]
  assign _T_565 = io_addr == 12'hb0f; // @[rvcsr.scala 380:61:@2231.4]
  assign _T_567 = io_addr == 12'hb8f; // @[rvcsr.scala 380:61:@2232.4]
  assign _T_569 = io_addr == 12'hb10; // @[rvcsr.scala 380:61:@2233.4]
  assign _T_571 = io_addr == 12'hb90; // @[rvcsr.scala 380:61:@2234.4]
  assign _T_573 = io_addr == 12'hb11; // @[rvcsr.scala 380:61:@2235.4]
  assign _T_575 = io_addr == 12'hb91; // @[rvcsr.scala 380:61:@2236.4]
  assign _T_577 = io_addr == 12'hb12; // @[rvcsr.scala 380:61:@2237.4]
  assign _T_579 = io_addr == 12'hb92; // @[rvcsr.scala 380:61:@2238.4]
  assign _T_581 = io_addr == 12'hb13; // @[rvcsr.scala 380:61:@2239.4]
  assign _T_583 = io_addr == 12'hb93; // @[rvcsr.scala 380:61:@2240.4]
  assign _T_585 = io_addr == 12'hb14; // @[rvcsr.scala 380:61:@2241.4]
  assign _T_587 = io_addr == 12'hb94; // @[rvcsr.scala 380:61:@2242.4]
  assign _T_589 = io_addr == 12'hb15; // @[rvcsr.scala 380:61:@2243.4]
  assign _T_591 = io_addr == 12'hb95; // @[rvcsr.scala 380:61:@2244.4]
  assign _T_593 = io_addr == 12'hb16; // @[rvcsr.scala 380:61:@2245.4]
  assign _T_595 = io_addr == 12'hb96; // @[rvcsr.scala 380:61:@2246.4]
  assign _T_597 = io_addr == 12'hb17; // @[rvcsr.scala 380:61:@2247.4]
  assign _T_599 = io_addr == 12'hb97; // @[rvcsr.scala 380:61:@2248.4]
  assign _T_601 = io_addr == 12'hb18; // @[rvcsr.scala 380:61:@2249.4]
  assign _T_603 = io_addr == 12'hb98; // @[rvcsr.scala 380:61:@2250.4]
  assign _T_605 = io_addr == 12'hb19; // @[rvcsr.scala 380:61:@2251.4]
  assign _T_607 = io_addr == 12'hb99; // @[rvcsr.scala 380:61:@2252.4]
  assign _T_609 = io_addr == 12'hb1a; // @[rvcsr.scala 380:61:@2253.4]
  assign _T_611 = io_addr == 12'hb9a; // @[rvcsr.scala 380:61:@2254.4]
  assign _T_613 = io_addr == 12'hb1b; // @[rvcsr.scala 380:61:@2255.4]
  assign _T_615 = io_addr == 12'hb9b; // @[rvcsr.scala 380:61:@2256.4]
  assign _T_617 = io_addr == 12'hb1c; // @[rvcsr.scala 380:61:@2257.4]
  assign _T_619 = io_addr == 12'hb9c; // @[rvcsr.scala 380:61:@2258.4]
  assign _T_621 = io_addr == 12'hb1d; // @[rvcsr.scala 380:61:@2259.4]
  assign _T_623 = io_addr == 12'hb9d; // @[rvcsr.scala 380:61:@2260.4]
  assign _T_625 = io_addr == 12'hb1e; // @[rvcsr.scala 380:61:@2261.4]
  assign _T_627 = io_addr == 12'hb9e; // @[rvcsr.scala 380:61:@2262.4]
  assign _T_629 = io_addr == 12'hb1f; // @[rvcsr.scala 380:61:@2263.4]
  assign _T_631 = io_addr == 12'hb9f; // @[rvcsr.scala 380:61:@2264.4]
  assign _T_633 = io_addr == 12'h323; // @[rvcsr.scala 380:61:@2265.4]
  assign _T_635 = io_addr == 12'h324; // @[rvcsr.scala 380:61:@2266.4]
  assign _T_637 = io_addr == 12'h325; // @[rvcsr.scala 380:61:@2267.4]
  assign _T_639 = io_addr == 12'h326; // @[rvcsr.scala 380:61:@2268.4]
  assign _T_641 = io_addr == 12'h327; // @[rvcsr.scala 380:61:@2269.4]
  assign _T_643 = io_addr == 12'h328; // @[rvcsr.scala 380:61:@2270.4]
  assign _T_645 = io_addr == 12'h329; // @[rvcsr.scala 380:61:@2271.4]
  assign _T_647 = io_addr == 12'h32a; // @[rvcsr.scala 380:61:@2272.4]
  assign _T_649 = io_addr == 12'h32b; // @[rvcsr.scala 380:61:@2273.4]
  assign _T_651 = io_addr == 12'h32c; // @[rvcsr.scala 380:61:@2274.4]
  assign _T_653 = io_addr == 12'h32d; // @[rvcsr.scala 380:61:@2275.4]
  assign _T_655 = io_addr == 12'h32e; // @[rvcsr.scala 380:61:@2276.4]
  assign _T_657 = io_addr == 12'h32f; // @[rvcsr.scala 380:61:@2277.4]
  assign _T_659 = io_addr == 12'h330; // @[rvcsr.scala 380:61:@2278.4]
  assign _T_661 = io_addr == 12'h331; // @[rvcsr.scala 380:61:@2279.4]
  assign _T_663 = io_addr == 12'h332; // @[rvcsr.scala 380:61:@2280.4]
  assign _T_665 = io_addr == 12'h333; // @[rvcsr.scala 380:61:@2281.4]
  assign _T_667 = io_addr == 12'h334; // @[rvcsr.scala 380:61:@2282.4]
  assign _T_669 = io_addr == 12'h335; // @[rvcsr.scala 380:61:@2283.4]
  assign _T_671 = io_addr == 12'h336; // @[rvcsr.scala 380:61:@2284.4]
  assign _T_673 = io_addr == 12'h337; // @[rvcsr.scala 380:61:@2285.4]
  assign _T_675 = io_addr == 12'h338; // @[rvcsr.scala 380:61:@2286.4]
  assign _T_677 = io_addr == 12'h339; // @[rvcsr.scala 380:61:@2287.4]
  assign _T_679 = io_addr == 12'h33a; // @[rvcsr.scala 380:61:@2288.4]
  assign _T_681 = io_addr == 12'h33b; // @[rvcsr.scala 380:61:@2289.4]
  assign _T_683 = io_addr == 12'h33c; // @[rvcsr.scala 380:61:@2290.4]
  assign _T_685 = io_addr == 12'h33d; // @[rvcsr.scala 380:61:@2291.4]
  assign _T_687 = io_addr == 12'h33e; // @[rvcsr.scala 380:61:@2292.4]
  assign _T_689 = io_addr == 12'h33f; // @[rvcsr.scala 380:61:@2293.4]
  assign _T_813 = 12'h33f == io_addr; // @[Mux.scala 46:19:@2302.4]
  assign _T_814 = _T_813 ? reg_mhpmevents_28 : 32'h0; // @[Mux.scala 46:16:@2303.4]
  assign _T_815 = 12'h33e == io_addr; // @[Mux.scala 46:19:@2304.4]
  assign _T_816 = _T_815 ? reg_mhpmevents_27 : _T_814; // @[Mux.scala 46:16:@2305.4]
  assign _T_817 = 12'h33d == io_addr; // @[Mux.scala 46:19:@2306.4]
  assign _T_818 = _T_817 ? reg_mhpmevents_26 : _T_816; // @[Mux.scala 46:16:@2307.4]
  assign _T_819 = 12'h33c == io_addr; // @[Mux.scala 46:19:@2308.4]
  assign _T_820 = _T_819 ? reg_mhpmevents_25 : _T_818; // @[Mux.scala 46:16:@2309.4]
  assign _T_821 = 12'h33b == io_addr; // @[Mux.scala 46:19:@2310.4]
  assign _T_822 = _T_821 ? reg_mhpmevents_24 : _T_820; // @[Mux.scala 46:16:@2311.4]
  assign _T_823 = 12'h33a == io_addr; // @[Mux.scala 46:19:@2312.4]
  assign _T_824 = _T_823 ? reg_mhpmevents_23 : _T_822; // @[Mux.scala 46:16:@2313.4]
  assign _T_825 = 12'h339 == io_addr; // @[Mux.scala 46:19:@2314.4]
  assign _T_826 = _T_825 ? reg_mhpmevents_22 : _T_824; // @[Mux.scala 46:16:@2315.4]
  assign _T_827 = 12'h338 == io_addr; // @[Mux.scala 46:19:@2316.4]
  assign _T_828 = _T_827 ? reg_mhpmevents_21 : _T_826; // @[Mux.scala 46:16:@2317.4]
  assign _T_829 = 12'h337 == io_addr; // @[Mux.scala 46:19:@2318.4]
  assign _T_830 = _T_829 ? reg_mhpmevents_20 : _T_828; // @[Mux.scala 46:16:@2319.4]
  assign _T_831 = 12'h336 == io_addr; // @[Mux.scala 46:19:@2320.4]
  assign _T_832 = _T_831 ? reg_mhpmevents_19 : _T_830; // @[Mux.scala 46:16:@2321.4]
  assign _T_833 = 12'h335 == io_addr; // @[Mux.scala 46:19:@2322.4]
  assign _T_834 = _T_833 ? reg_mhpmevents_18 : _T_832; // @[Mux.scala 46:16:@2323.4]
  assign _T_835 = 12'h334 == io_addr; // @[Mux.scala 46:19:@2324.4]
  assign _T_836 = _T_835 ? reg_mhpmevents_17 : _T_834; // @[Mux.scala 46:16:@2325.4]
  assign _T_837 = 12'h333 == io_addr; // @[Mux.scala 46:19:@2326.4]
  assign _T_838 = _T_837 ? reg_mhpmevents_16 : _T_836; // @[Mux.scala 46:16:@2327.4]
  assign _T_839 = 12'h332 == io_addr; // @[Mux.scala 46:19:@2328.4]
  assign _T_840 = _T_839 ? reg_mhpmevents_15 : _T_838; // @[Mux.scala 46:16:@2329.4]
  assign _T_841 = 12'h331 == io_addr; // @[Mux.scala 46:19:@2330.4]
  assign _T_842 = _T_841 ? reg_mhpmevents_14 : _T_840; // @[Mux.scala 46:16:@2331.4]
  assign _T_843 = 12'h330 == io_addr; // @[Mux.scala 46:19:@2332.4]
  assign _T_844 = _T_843 ? reg_mhpmevents_13 : _T_842; // @[Mux.scala 46:16:@2333.4]
  assign _T_845 = 12'h32f == io_addr; // @[Mux.scala 46:19:@2334.4]
  assign _T_846 = _T_845 ? reg_mhpmevents_12 : _T_844; // @[Mux.scala 46:16:@2335.4]
  assign _T_847 = 12'h32e == io_addr; // @[Mux.scala 46:19:@2336.4]
  assign _T_848 = _T_847 ? reg_mhpmevents_11 : _T_846; // @[Mux.scala 46:16:@2337.4]
  assign _T_849 = 12'h32d == io_addr; // @[Mux.scala 46:19:@2338.4]
  assign _T_850 = _T_849 ? reg_mhpmevents_10 : _T_848; // @[Mux.scala 46:16:@2339.4]
  assign _T_851 = 12'h32c == io_addr; // @[Mux.scala 46:19:@2340.4]
  assign _T_852 = _T_851 ? reg_mhpmevents_9 : _T_850; // @[Mux.scala 46:16:@2341.4]
  assign _T_853 = 12'h32b == io_addr; // @[Mux.scala 46:19:@2342.4]
  assign _T_854 = _T_853 ? reg_mhpmevents_8 : _T_852; // @[Mux.scala 46:16:@2343.4]
  assign _T_855 = 12'h32a == io_addr; // @[Mux.scala 46:19:@2344.4]
  assign _T_856 = _T_855 ? reg_mhpmevents_7 : _T_854; // @[Mux.scala 46:16:@2345.4]
  assign _T_857 = 12'h329 == io_addr; // @[Mux.scala 46:19:@2346.4]
  assign _T_858 = _T_857 ? reg_mhpmevents_6 : _T_856; // @[Mux.scala 46:16:@2347.4]
  assign _T_859 = 12'h328 == io_addr; // @[Mux.scala 46:19:@2348.4]
  assign _T_860 = _T_859 ? reg_mhpmevents_5 : _T_858; // @[Mux.scala 46:16:@2349.4]
  assign _T_861 = 12'h327 == io_addr; // @[Mux.scala 46:19:@2350.4]
  assign _T_862 = _T_861 ? reg_mhpmevents_4 : _T_860; // @[Mux.scala 46:16:@2351.4]
  assign _T_863 = 12'h326 == io_addr; // @[Mux.scala 46:19:@2352.4]
  assign _T_864 = _T_863 ? reg_mhpmevents_3 : _T_862; // @[Mux.scala 46:16:@2353.4]
  assign _T_865 = 12'h325 == io_addr; // @[Mux.scala 46:19:@2354.4]
  assign _T_866 = _T_865 ? reg_mhpmevents_2 : _T_864; // @[Mux.scala 46:16:@2355.4]
  assign _T_867 = 12'h324 == io_addr; // @[Mux.scala 46:19:@2356.4]
  assign _T_868 = _T_867 ? reg_mhpmevents_1 : _T_866; // @[Mux.scala 46:16:@2357.4]
  assign _T_869 = 12'h323 == io_addr; // @[Mux.scala 46:19:@2358.4]
  assign _T_870 = _T_869 ? reg_mhpmevents_0 : _T_868; // @[Mux.scala 46:16:@2359.4]
  assign _T_871 = 12'hb9f == io_addr; // @[Mux.scala 46:19:@2360.4]
  assign _T_872 = _T_871 ? _T_172 : _T_870; // @[Mux.scala 46:16:@2361.4]
  assign _T_873 = 12'hb1f == io_addr; // @[Mux.scala 46:19:@2362.4]
  assign _T_874 = _T_873 ? _T_171 : _T_872; // @[Mux.scala 46:16:@2363.4]
  assign _T_875 = 12'hb9e == io_addr; // @[Mux.scala 46:19:@2364.4]
  assign _T_876 = _T_875 ? _T_170 : _T_874; // @[Mux.scala 46:16:@2365.4]
  assign _T_877 = 12'hb1e == io_addr; // @[Mux.scala 46:19:@2366.4]
  assign _T_878 = _T_877 ? _T_169 : _T_876; // @[Mux.scala 46:16:@2367.4]
  assign _T_879 = 12'hb9d == io_addr; // @[Mux.scala 46:19:@2368.4]
  assign _T_880 = _T_879 ? _T_168 : _T_878; // @[Mux.scala 46:16:@2369.4]
  assign _T_881 = 12'hb1d == io_addr; // @[Mux.scala 46:19:@2370.4]
  assign _T_882 = _T_881 ? _T_167 : _T_880; // @[Mux.scala 46:16:@2371.4]
  assign _T_883 = 12'hb9c == io_addr; // @[Mux.scala 46:19:@2372.4]
  assign _T_884 = _T_883 ? _T_166 : _T_882; // @[Mux.scala 46:16:@2373.4]
  assign _T_885 = 12'hb1c == io_addr; // @[Mux.scala 46:19:@2374.4]
  assign _T_886 = _T_885 ? _T_165 : _T_884; // @[Mux.scala 46:16:@2375.4]
  assign _T_887 = 12'hb9b == io_addr; // @[Mux.scala 46:19:@2376.4]
  assign _T_888 = _T_887 ? _T_164 : _T_886; // @[Mux.scala 46:16:@2377.4]
  assign _T_889 = 12'hb1b == io_addr; // @[Mux.scala 46:19:@2378.4]
  assign _T_890 = _T_889 ? _T_163 : _T_888; // @[Mux.scala 46:16:@2379.4]
  assign _T_891 = 12'hb9a == io_addr; // @[Mux.scala 46:19:@2380.4]
  assign _T_892 = _T_891 ? _T_162 : _T_890; // @[Mux.scala 46:16:@2381.4]
  assign _T_893 = 12'hb1a == io_addr; // @[Mux.scala 46:19:@2382.4]
  assign _T_894 = _T_893 ? _T_161 : _T_892; // @[Mux.scala 46:16:@2383.4]
  assign _T_895 = 12'hb99 == io_addr; // @[Mux.scala 46:19:@2384.4]
  assign _T_896 = _T_895 ? _T_160 : _T_894; // @[Mux.scala 46:16:@2385.4]
  assign _T_897 = 12'hb19 == io_addr; // @[Mux.scala 46:19:@2386.4]
  assign _T_898 = _T_897 ? _T_159 : _T_896; // @[Mux.scala 46:16:@2387.4]
  assign _T_899 = 12'hb98 == io_addr; // @[Mux.scala 46:19:@2388.4]
  assign _T_900 = _T_899 ? _T_158 : _T_898; // @[Mux.scala 46:16:@2389.4]
  assign _T_901 = 12'hb18 == io_addr; // @[Mux.scala 46:19:@2390.4]
  assign _T_902 = _T_901 ? _T_157 : _T_900; // @[Mux.scala 46:16:@2391.4]
  assign _T_903 = 12'hb97 == io_addr; // @[Mux.scala 46:19:@2392.4]
  assign _T_904 = _T_903 ? _T_156 : _T_902; // @[Mux.scala 46:16:@2393.4]
  assign _T_905 = 12'hb17 == io_addr; // @[Mux.scala 46:19:@2394.4]
  assign _T_906 = _T_905 ? _T_155 : _T_904; // @[Mux.scala 46:16:@2395.4]
  assign _T_907 = 12'hb96 == io_addr; // @[Mux.scala 46:19:@2396.4]
  assign _T_908 = _T_907 ? _T_154 : _T_906; // @[Mux.scala 46:16:@2397.4]
  assign _T_909 = 12'hb16 == io_addr; // @[Mux.scala 46:19:@2398.4]
  assign _T_910 = _T_909 ? _T_153 : _T_908; // @[Mux.scala 46:16:@2399.4]
  assign _T_911 = 12'hb95 == io_addr; // @[Mux.scala 46:19:@2400.4]
  assign _T_912 = _T_911 ? _T_152 : _T_910; // @[Mux.scala 46:16:@2401.4]
  assign _T_913 = 12'hb15 == io_addr; // @[Mux.scala 46:19:@2402.4]
  assign _T_914 = _T_913 ? _T_151 : _T_912; // @[Mux.scala 46:16:@2403.4]
  assign _T_915 = 12'hb94 == io_addr; // @[Mux.scala 46:19:@2404.4]
  assign _T_916 = _T_915 ? _T_150 : _T_914; // @[Mux.scala 46:16:@2405.4]
  assign _T_917 = 12'hb14 == io_addr; // @[Mux.scala 46:19:@2406.4]
  assign _T_918 = _T_917 ? _T_149 : _T_916; // @[Mux.scala 46:16:@2407.4]
  assign _T_919 = 12'hb93 == io_addr; // @[Mux.scala 46:19:@2408.4]
  assign _T_920 = _T_919 ? _T_148 : _T_918; // @[Mux.scala 46:16:@2409.4]
  assign _T_921 = 12'hb13 == io_addr; // @[Mux.scala 46:19:@2410.4]
  assign _T_922 = _T_921 ? _T_147 : _T_920; // @[Mux.scala 46:16:@2411.4]
  assign _T_923 = 12'hb92 == io_addr; // @[Mux.scala 46:19:@2412.4]
  assign _T_924 = _T_923 ? _T_146 : _T_922; // @[Mux.scala 46:16:@2413.4]
  assign _T_925 = 12'hb12 == io_addr; // @[Mux.scala 46:19:@2414.4]
  assign _T_926 = _T_925 ? _T_145 : _T_924; // @[Mux.scala 46:16:@2415.4]
  assign _T_927 = 12'hb91 == io_addr; // @[Mux.scala 46:19:@2416.4]
  assign _T_928 = _T_927 ? _T_144 : _T_926; // @[Mux.scala 46:16:@2417.4]
  assign _T_929 = 12'hb11 == io_addr; // @[Mux.scala 46:19:@2418.4]
  assign _T_930 = _T_929 ? _T_143 : _T_928; // @[Mux.scala 46:16:@2419.4]
  assign _T_931 = 12'hb90 == io_addr; // @[Mux.scala 46:19:@2420.4]
  assign _T_932 = _T_931 ? _T_142 : _T_930; // @[Mux.scala 46:16:@2421.4]
  assign _T_933 = 12'hb10 == io_addr; // @[Mux.scala 46:19:@2422.4]
  assign _T_934 = _T_933 ? _T_141 : _T_932; // @[Mux.scala 46:16:@2423.4]
  assign _T_935 = 12'hb8f == io_addr; // @[Mux.scala 46:19:@2424.4]
  assign _T_936 = _T_935 ? _T_140 : _T_934; // @[Mux.scala 46:16:@2425.4]
  assign _T_937 = 12'hb0f == io_addr; // @[Mux.scala 46:19:@2426.4]
  assign _T_938 = _T_937 ? _T_139 : _T_936; // @[Mux.scala 46:16:@2427.4]
  assign _T_939 = 12'hb8e == io_addr; // @[Mux.scala 46:19:@2428.4]
  assign _T_940 = _T_939 ? _T_138 : _T_938; // @[Mux.scala 46:16:@2429.4]
  assign _T_941 = 12'hb0e == io_addr; // @[Mux.scala 46:19:@2430.4]
  assign _T_942 = _T_941 ? _T_137 : _T_940; // @[Mux.scala 46:16:@2431.4]
  assign _T_943 = 12'hb8d == io_addr; // @[Mux.scala 46:19:@2432.4]
  assign _T_944 = _T_943 ? _T_136 : _T_942; // @[Mux.scala 46:16:@2433.4]
  assign _T_945 = 12'hb0d == io_addr; // @[Mux.scala 46:19:@2434.4]
  assign _T_946 = _T_945 ? _T_135 : _T_944; // @[Mux.scala 46:16:@2435.4]
  assign _T_947 = 12'hb8c == io_addr; // @[Mux.scala 46:19:@2436.4]
  assign _T_948 = _T_947 ? _T_134 : _T_946; // @[Mux.scala 46:16:@2437.4]
  assign _T_949 = 12'hb0c == io_addr; // @[Mux.scala 46:19:@2438.4]
  assign _T_950 = _T_949 ? _T_133 : _T_948; // @[Mux.scala 46:16:@2439.4]
  assign _T_951 = 12'hb8b == io_addr; // @[Mux.scala 46:19:@2440.4]
  assign _T_952 = _T_951 ? _T_132 : _T_950; // @[Mux.scala 46:16:@2441.4]
  assign _T_953 = 12'hb0b == io_addr; // @[Mux.scala 46:19:@2442.4]
  assign _T_954 = _T_953 ? _T_131 : _T_952; // @[Mux.scala 46:16:@2443.4]
  assign _T_955 = 12'hb8a == io_addr; // @[Mux.scala 46:19:@2444.4]
  assign _T_956 = _T_955 ? _T_130 : _T_954; // @[Mux.scala 46:16:@2445.4]
  assign _T_957 = 12'hb0a == io_addr; // @[Mux.scala 46:19:@2446.4]
  assign _T_958 = _T_957 ? _T_129 : _T_956; // @[Mux.scala 46:16:@2447.4]
  assign _T_959 = 12'hb89 == io_addr; // @[Mux.scala 46:19:@2448.4]
  assign _T_960 = _T_959 ? _T_128 : _T_958; // @[Mux.scala 46:16:@2449.4]
  assign _T_961 = 12'hb09 == io_addr; // @[Mux.scala 46:19:@2450.4]
  assign _T_962 = _T_961 ? _T_127 : _T_960; // @[Mux.scala 46:16:@2451.4]
  assign _T_963 = 12'hb88 == io_addr; // @[Mux.scala 46:19:@2452.4]
  assign _T_964 = _T_963 ? _T_126 : _T_962; // @[Mux.scala 46:16:@2453.4]
  assign _T_965 = 12'hb08 == io_addr; // @[Mux.scala 46:19:@2454.4]
  assign _T_966 = _T_965 ? _T_125 : _T_964; // @[Mux.scala 46:16:@2455.4]
  assign _T_967 = 12'hb87 == io_addr; // @[Mux.scala 46:19:@2456.4]
  assign _T_968 = _T_967 ? _T_124 : _T_966; // @[Mux.scala 46:16:@2457.4]
  assign _T_969 = 12'hb07 == io_addr; // @[Mux.scala 46:19:@2458.4]
  assign _T_970 = _T_969 ? _T_123 : _T_968; // @[Mux.scala 46:16:@2459.4]
  assign _T_971 = 12'hb86 == io_addr; // @[Mux.scala 46:19:@2460.4]
  assign _T_972 = _T_971 ? _T_122 : _T_970; // @[Mux.scala 46:16:@2461.4]
  assign _T_973 = 12'hb06 == io_addr; // @[Mux.scala 46:19:@2462.4]
  assign _T_974 = _T_973 ? _T_121 : _T_972; // @[Mux.scala 46:16:@2463.4]
  assign _T_975 = 12'hb85 == io_addr; // @[Mux.scala 46:19:@2464.4]
  assign _T_976 = _T_975 ? _T_120 : _T_974; // @[Mux.scala 46:16:@2465.4]
  assign _T_977 = 12'hb05 == io_addr; // @[Mux.scala 46:19:@2466.4]
  assign _T_978 = _T_977 ? _T_119 : _T_976; // @[Mux.scala 46:16:@2467.4]
  assign _T_979 = 12'hb84 == io_addr; // @[Mux.scala 46:19:@2468.4]
  assign _T_980 = _T_979 ? _T_118 : _T_978; // @[Mux.scala 46:16:@2469.4]
  assign _T_981 = 12'hb04 == io_addr; // @[Mux.scala 46:19:@2470.4]
  assign _T_982 = _T_981 ? _T_117 : _T_980; // @[Mux.scala 46:16:@2471.4]
  assign _T_983 = 12'hb83 == io_addr; // @[Mux.scala 46:19:@2472.4]
  assign _T_984 = _T_983 ? _T_116 : _T_982; // @[Mux.scala 46:16:@2473.4]
  assign _T_985 = 12'hb03 == io_addr; // @[Mux.scala 46:19:@2474.4]
  assign _T_986 = _T_985 ? _T_115 : _T_984; // @[Mux.scala 46:16:@2475.4]
  assign _T_987 = 12'h7b3 == io_addr; // @[Mux.scala 46:19:@2476.4]
  assign _T_988 = _T_987 ? reg_dscratch1 : _T_986; // @[Mux.scala 46:16:@2477.4]
  assign _T_989 = 12'h7b2 == io_addr; // @[Mux.scala 46:19:@2478.4]
  assign _T_990 = _T_989 ? reg_dscratch0 : _T_988; // @[Mux.scala 46:16:@2479.4]
  assign _T_991 = 12'h7b1 == io_addr; // @[Mux.scala 46:19:@2480.4]
  assign _T_992 = _T_991 ? reg_dpc : _T_990; // @[Mux.scala 46:16:@2481.4]
  assign _T_993 = 12'h7b0 == io_addr; // @[Mux.scala 46:19:@2482.4]
  assign _T_994 = _T_993 ? reg_dcsr : _T_992; // @[Mux.scala 46:16:@2483.4]
  assign _T_995 = 12'hba0 == io_addr; // @[Mux.scala 46:19:@2484.4]
  assign _T_996 = _T_995 ? _T_112 : _T_994; // @[Mux.scala 46:16:@2485.4]
  assign _T_997 = 12'hb81 == io_addr; // @[Mux.scala 46:19:@2486.4]
  assign _T_998 = _T_997 ? _T_113 : _T_996; // @[Mux.scala 46:16:@2487.4]
  assign _T_999 = 12'hb20 == io_addr; // @[Mux.scala 46:19:@2488.4]
  assign _T_1000 = _T_999 ? _T_112 : _T_998; // @[Mux.scala 46:16:@2489.4]
  assign _T_1001 = 12'hb01 == io_addr; // @[Mux.scala 46:19:@2490.4]
  assign _T_1002 = _T_1001 ? _T_111 : _T_1000; // @[Mux.scala 46:16:@2491.4]
  assign _T_1003 = 12'hb82 == io_addr; // @[Mux.scala 46:19:@2492.4]
  assign _T_1004 = _T_1003 ? _T_108 : _T_1002; // @[Mux.scala 46:16:@2493.4]
  assign _T_1005 = 12'hb80 == io_addr; // @[Mux.scala 46:19:@2494.4]
  assign _T_1006 = _T_1005 ? _T_107 : _T_1004; // @[Mux.scala 46:16:@2495.4]
  assign _T_1007 = 12'hb02 == io_addr; // @[Mux.scala 46:19:@2496.4]
  assign _T_1008 = _T_1007 ? _T_108 : _T_1006; // @[Mux.scala 46:16:@2497.4]
  assign _T_1009 = 12'hb00 == io_addr; // @[Mux.scala 46:19:@2498.4]
  assign _T_1010 = _T_1009 ? _T_107 : _T_1008; // @[Mux.scala 46:16:@2499.4]
  assign _T_1011 = 12'h344 == io_addr; // @[Mux.scala 46:19:@2500.4]
  assign _T_1012 = _T_1011 ? reg_mip : _T_1010; // @[Mux.scala 46:16:@2501.4]
  assign _T_1013 = 12'h343 == io_addr; // @[Mux.scala 46:19:@2502.4]
  assign _T_1014 = _T_1013 ? reg_mtval : _T_1012; // @[Mux.scala 46:16:@2503.4]
  assign _T_1015 = 12'h342 == io_addr; // @[Mux.scala 46:19:@2504.4]
  assign _T_1016 = _T_1015 ? reg_mcause : _T_1014; // @[Mux.scala 46:16:@2505.4]
  assign _T_1017 = 12'h341 == io_addr; // @[Mux.scala 46:19:@2506.4]
  assign _T_1018 = _T_1017 ? reg_mepc : _T_1016; // @[Mux.scala 46:16:@2507.4]
  assign _T_1019 = 12'h340 == io_addr; // @[Mux.scala 46:19:@2508.4]
  assign _T_1020 = _T_1019 ? reg_mscratch : _T_1018; // @[Mux.scala 46:16:@2509.4]
  assign _T_1021 = 12'h306 == io_addr; // @[Mux.scala 46:19:@2510.4]
  assign _T_1022 = _T_1021 ? reg_mcounteren : _T_1020; // @[Mux.scala 46:16:@2511.4]
  assign _T_1023 = 12'h305 == io_addr; // @[Mux.scala 46:19:@2512.4]
  assign _T_1024 = _T_1023 ? reg_mtvec : _T_1022; // @[Mux.scala 46:16:@2513.4]
  assign _T_1025 = 12'h304 == io_addr; // @[Mux.scala 46:19:@2514.4]
  assign _T_1026 = _T_1025 ? reg_mie : _T_1024; // @[Mux.scala 46:16:@2515.4]
  assign _T_1027 = 12'h303 == io_addr; // @[Mux.scala 46:19:@2516.4]
  assign _T_1028 = _T_1027 ? reg_mideleg : _T_1026; // @[Mux.scala 46:16:@2517.4]
  assign _T_1029 = 12'h302 == io_addr; // @[Mux.scala 46:19:@2518.4]
  assign _T_1030 = _T_1029 ? reg_medeleg : _T_1028; // @[Mux.scala 46:16:@2519.4]
  assign _T_1031 = 12'h301 == io_addr; // @[Mux.scala 46:19:@2520.4]
  assign _T_1032 = _T_1031 ? 32'h40000100 : _T_1030; // @[Mux.scala 46:16:@2521.4]
  assign _T_1033 = 12'h300 == io_addr; // @[Mux.scala 46:19:@2522.4]
  assign _T_1034 = _T_1033 ? reg_mstatus : _T_1032; // @[Mux.scala 46:16:@2523.4]
  assign _T_1035 = 12'hf14 == io_addr; // @[Mux.scala 46:19:@2524.4]
  assign _T_1036 = _T_1035 ? 32'h0 : _T_1034; // @[Mux.scala 46:16:@2525.4]
  assign _T_1037 = 12'hf13 == io_addr; // @[Mux.scala 46:19:@2526.4]
  assign _T_1038 = _T_1037 ? 32'h8000 : _T_1036; // @[Mux.scala 46:16:@2527.4]
  assign _T_1039 = 12'hf12 == io_addr; // @[Mux.scala 46:19:@2528.4]
  assign _T_1040 = _T_1039 ? 32'h0 : _T_1038; // @[Mux.scala 46:16:@2529.4]
  assign _T_1041 = 12'hf11 == io_addr; // @[Mux.scala 46:19:@2530.4]
  assign _T_1042 = _T_1041 ? 32'h0 : _T_1040; // @[Mux.scala 46:16:@2531.4]
  assign _T_1044 = legal_priv ? _T_1042 : 32'h0; // @[rvcsr.scala 389:20:@2532.4]
  assign _T_1065 = csr_wdata[2]; // @[rvcsr.scala 396:55:@2554.8]
  assign _GEN_56 = _T_469 ? _T_447 : _GEN_38; // @[rvcsr.scala 395:41:@2546.6]
  assign _T_1122 = {mie_rsrvd4,mie_SSIE}; // @[rvcsr.scala 407:28:@2648.8]
  assign _T_1123 = {_T_1122,mie_USIE}; // @[rvcsr.scala 407:28:@2649.8]
  assign _T_1124 = {mie_STIE,mie_UTIE}; // @[rvcsr.scala 407:28:@2650.8]
  assign _GEN_58 = _T_477 ? _T_1156 : _T_348; // @[rvcsr.scala 402:37:@2616.6]
  assign mie_MSIE = csr_wen ? _GEN_58 : _T_348; // @[rvcsr.scala 393:19:@2545.4]
  assign _T_1125 = {_T_1124,mie_MSIE}; // @[rvcsr.scala 407:28:@2651.8]
  assign _T_1126 = {_T_1125,_T_1123}; // @[rvcsr.scala 407:28:@2652.8]
  assign _GEN_57 = _T_477 ? _T_1160 : _T_352; // @[rvcsr.scala 402:37:@2616.6]
  assign mie_MTIE = csr_wen ? _GEN_57 : _T_352; // @[rvcsr.scala 393:19:@2545.4]
  assign _T_1127 = {mie_UEIE,mie_MTIE}; // @[rvcsr.scala 407:28:@2653.8]
  assign _T_1128 = {_T_1127,mie_rsrvd3}; // @[rvcsr.scala 407:28:@2654.8]
  assign _T_1129 = {mie_rsrvd2,mie_SEIE}; // @[rvcsr.scala 407:28:@2655.8]
  assign _T_1130 = {mie_rsrvd1,mie_MEIE}; // @[rvcsr.scala 407:28:@2656.8]
  assign _T_1131 = {_T_1130,_T_1129}; // @[rvcsr.scala 407:28:@2657.8]
  assign _T_1132 = {_T_1131,_T_1128}; // @[rvcsr.scala 407:28:@2658.8]
  assign _T_1133 = {_T_1132,_T_1126}; // @[rvcsr.scala 407:28:@2659.8]
  assign _GEN_59 = _T_477 ? {{1'd0}, _T_1133} : reg_mie; // @[rvcsr.scala 402:37:@2616.6]
  assign _T_1134 = csr_wdata[31:2]; // @[rvcsr.scala 411:39:@2663.8]
  assign _T_1140 = {_T_1134,2'h0}; // @[Cat.scala 30:58:@2665.8]
  assign _GEN_60 = _T_479 ? _T_1140 : reg_mtvec; // @[rvcsr.scala 410:39:@2662.6]
  assign _GEN_61 = _T_481 ? csr_wdata : reg_mcounteren; // @[rvcsr.scala 414:44:@2668.6]
  assign _GEN_62 = _T_483 ? csr_wdata : reg_mscratch; // @[rvcsr.scala 418:42:@2671.6]
  assign _GEN_63 = _T_485 ? _T_1140 : _GEN_52; // @[rvcsr.scala 422:38:@2674.6]
  assign _GEN_64 = _T_487 ? csr_wdata : _GEN_51; // @[rvcsr.scala 426:40:@2680.6]
  assign _GEN_65 = _T_489 ? csr_wdata : reg_mtval; // @[rvcsr.scala 430:39:@2683.6]
  assign _GEN_68 = _T_491 ? {{1'd0}, _T_420} : _GEN_33; // @[rvcsr.scala 434:37:@2686.6]
  assign _T_1178 = reg_mcycle[63:32]; // @[rvcsr.scala 444:41:@2733.8]
  assign _T_1179 = {_T_1178,csr_wdata}; // @[Cat.scala 30:58:@2734.8]
  assign _GEN_69 = _T_493 ? _T_1179 : _GEN_0; // @[rvcsr.scala 442:40:@2732.6]
  assign _T_1181 = {_T_108,csr_wdata}; // @[Cat.scala 30:58:@2739.8]
  assign _GEN_70 = _T_495 ? _T_1181 : _GEN_2; // @[rvcsr.scala 447:42:@2737.6]
  assign _T_1183 = {csr_wdata,_T_107}; // @[Cat.scala 30:58:@2744.8]
  assign _GEN_71 = _T_497 ? _T_1183 : _GEN_69; // @[rvcsr.scala 452:41:@2742.6]
  assign _T_1184 = reg_minstret[31:0]; // @[rvcsr.scala 459:56:@2748.8]
  assign _T_1185 = {csr_wdata,_T_1184}; // @[Cat.scala 30:58:@2749.8]
  assign _GEN_72 = _T_499 ? _T_1185 : _GEN_70; // @[rvcsr.scala 457:43:@2747.6]
  assign _T_1187 = {_T_116,csr_wdata}; // @[Cat.scala 30:58:@2754.8]
  assign _GEN_73 = _T_517 ? _T_1187 : _GEN_3; // @[rvcsr.scala 463:57:@2752.6]
  assign _T_1189 = {_T_118,csr_wdata}; // @[Cat.scala 30:58:@2759.8]
  assign _GEN_74 = _T_521 ? _T_1189 : _GEN_4; // @[rvcsr.scala 463:57:@2757.6]
  assign _T_1191 = {_T_120,csr_wdata}; // @[Cat.scala 30:58:@2764.8]
  assign _GEN_75 = _T_525 ? _T_1191 : _GEN_5; // @[rvcsr.scala 463:57:@2762.6]
  assign _T_1193 = {_T_122,csr_wdata}; // @[Cat.scala 30:58:@2769.8]
  assign _GEN_76 = _T_529 ? _T_1193 : _GEN_6; // @[rvcsr.scala 463:57:@2767.6]
  assign _T_1195 = {_T_124,csr_wdata}; // @[Cat.scala 30:58:@2774.8]
  assign _GEN_77 = _T_533 ? _T_1195 : _GEN_7; // @[rvcsr.scala 463:57:@2772.6]
  assign _T_1197 = {_T_126,csr_wdata}; // @[Cat.scala 30:58:@2779.8]
  assign _GEN_78 = _T_537 ? _T_1197 : _GEN_8; // @[rvcsr.scala 463:57:@2777.6]
  assign _T_1199 = {_T_128,csr_wdata}; // @[Cat.scala 30:58:@2784.8]
  assign _GEN_79 = _T_541 ? _T_1199 : _GEN_9; // @[rvcsr.scala 463:57:@2782.6]
  assign _T_1201 = {_T_130,csr_wdata}; // @[Cat.scala 30:58:@2789.8]
  assign _GEN_80 = _T_545 ? _T_1201 : _GEN_10; // @[rvcsr.scala 463:57:@2787.6]
  assign _T_1203 = {_T_132,csr_wdata}; // @[Cat.scala 30:58:@2794.8]
  assign _GEN_81 = _T_549 ? _T_1203 : _GEN_11; // @[rvcsr.scala 463:57:@2792.6]
  assign _T_1205 = {_T_134,csr_wdata}; // @[Cat.scala 30:58:@2799.8]
  assign _GEN_82 = _T_553 ? _T_1205 : _GEN_12; // @[rvcsr.scala 463:57:@2797.6]
  assign _T_1207 = {_T_136,csr_wdata}; // @[Cat.scala 30:58:@2804.8]
  assign _GEN_83 = _T_557 ? _T_1207 : _GEN_13; // @[rvcsr.scala 463:57:@2802.6]
  assign _T_1209 = {_T_138,csr_wdata}; // @[Cat.scala 30:58:@2809.8]
  assign _GEN_84 = _T_561 ? _T_1209 : _GEN_14; // @[rvcsr.scala 463:57:@2807.6]
  assign _T_1211 = {_T_140,csr_wdata}; // @[Cat.scala 30:58:@2814.8]
  assign _GEN_85 = _T_565 ? _T_1211 : _GEN_15; // @[rvcsr.scala 463:57:@2812.6]
  assign _T_1213 = {_T_142,csr_wdata}; // @[Cat.scala 30:58:@2819.8]
  assign _GEN_86 = _T_569 ? _T_1213 : _GEN_16; // @[rvcsr.scala 463:57:@2817.6]
  assign _T_1215 = {_T_144,csr_wdata}; // @[Cat.scala 30:58:@2824.8]
  assign _GEN_87 = _T_573 ? _T_1215 : _GEN_17; // @[rvcsr.scala 463:57:@2822.6]
  assign _T_1217 = {_T_146,csr_wdata}; // @[Cat.scala 30:58:@2829.8]
  assign _GEN_88 = _T_577 ? _T_1217 : _GEN_18; // @[rvcsr.scala 463:57:@2827.6]
  assign _T_1219 = {_T_148,csr_wdata}; // @[Cat.scala 30:58:@2834.8]
  assign _GEN_89 = _T_581 ? _T_1219 : _GEN_19; // @[rvcsr.scala 463:57:@2832.6]
  assign _T_1221 = {_T_150,csr_wdata}; // @[Cat.scala 30:58:@2839.8]
  assign _GEN_90 = _T_585 ? _T_1221 : _GEN_20; // @[rvcsr.scala 463:57:@2837.6]
  assign _T_1223 = {_T_152,csr_wdata}; // @[Cat.scala 30:58:@2844.8]
  assign _GEN_91 = _T_589 ? _T_1223 : _GEN_21; // @[rvcsr.scala 463:57:@2842.6]
  assign _T_1225 = {_T_154,csr_wdata}; // @[Cat.scala 30:58:@2849.8]
  assign _GEN_92 = _T_593 ? _T_1225 : _GEN_22; // @[rvcsr.scala 463:57:@2847.6]
  assign _T_1227 = {_T_156,csr_wdata}; // @[Cat.scala 30:58:@2854.8]
  assign _GEN_93 = _T_597 ? _T_1227 : _GEN_23; // @[rvcsr.scala 463:57:@2852.6]
  assign _T_1229 = {_T_158,csr_wdata}; // @[Cat.scala 30:58:@2859.8]
  assign _GEN_94 = _T_601 ? _T_1229 : _GEN_24; // @[rvcsr.scala 463:57:@2857.6]
  assign _T_1231 = {_T_160,csr_wdata}; // @[Cat.scala 30:58:@2864.8]
  assign _GEN_95 = _T_605 ? _T_1231 : _GEN_25; // @[rvcsr.scala 463:57:@2862.6]
  assign _T_1233 = {_T_162,csr_wdata}; // @[Cat.scala 30:58:@2869.8]
  assign _GEN_96 = _T_609 ? _T_1233 : _GEN_26; // @[rvcsr.scala 463:57:@2867.6]
  assign _T_1235 = {_T_164,csr_wdata}; // @[Cat.scala 30:58:@2874.8]
  assign _GEN_97 = _T_613 ? _T_1235 : _GEN_27; // @[rvcsr.scala 463:57:@2872.6]
  assign _T_1237 = {_T_166,csr_wdata}; // @[Cat.scala 30:58:@2879.8]
  assign _GEN_98 = _T_617 ? _T_1237 : _GEN_28; // @[rvcsr.scala 463:57:@2877.6]
  assign _T_1239 = {_T_168,csr_wdata}; // @[Cat.scala 30:58:@2884.8]
  assign _GEN_99 = _T_621 ? _T_1239 : _GEN_29; // @[rvcsr.scala 463:57:@2882.6]
  assign _T_1241 = {_T_170,csr_wdata}; // @[Cat.scala 30:58:@2889.8]
  assign _GEN_100 = _T_625 ? _T_1241 : _GEN_30; // @[rvcsr.scala 463:57:@2887.6]
  assign _T_1243 = {_T_172,csr_wdata}; // @[Cat.scala 30:58:@2894.8]
  assign _GEN_101 = _T_629 ? _T_1243 : _GEN_31; // @[rvcsr.scala 463:57:@2892.6]
  assign _T_1245 = {csr_wdata,_T_115}; // @[Cat.scala 30:58:@2899.8]
  assign _GEN_102 = _T_519 ? _T_1245 : _GEN_73; // @[rvcsr.scala 470:58:@2897.6]
  assign _T_1247 = {csr_wdata,_T_117}; // @[Cat.scala 30:58:@2904.8]
  assign _GEN_103 = _T_523 ? _T_1247 : _GEN_74; // @[rvcsr.scala 470:58:@2902.6]
  assign _T_1249 = {csr_wdata,_T_119}; // @[Cat.scala 30:58:@2909.8]
  assign _GEN_104 = _T_527 ? _T_1249 : _GEN_75; // @[rvcsr.scala 470:58:@2907.6]
  assign _T_1251 = {csr_wdata,_T_121}; // @[Cat.scala 30:58:@2914.8]
  assign _GEN_105 = _T_531 ? _T_1251 : _GEN_76; // @[rvcsr.scala 470:58:@2912.6]
  assign _T_1253 = {csr_wdata,_T_123}; // @[Cat.scala 30:58:@2919.8]
  assign _GEN_106 = _T_535 ? _T_1253 : _GEN_77; // @[rvcsr.scala 470:58:@2917.6]
  assign _T_1255 = {csr_wdata,_T_125}; // @[Cat.scala 30:58:@2924.8]
  assign _GEN_107 = _T_539 ? _T_1255 : _GEN_78; // @[rvcsr.scala 470:58:@2922.6]
  assign _T_1257 = {csr_wdata,_T_127}; // @[Cat.scala 30:58:@2929.8]
  assign _GEN_108 = _T_543 ? _T_1257 : _GEN_79; // @[rvcsr.scala 470:58:@2927.6]
  assign _T_1259 = {csr_wdata,_T_129}; // @[Cat.scala 30:58:@2934.8]
  assign _GEN_109 = _T_547 ? _T_1259 : _GEN_80; // @[rvcsr.scala 470:58:@2932.6]
  assign _T_1261 = {csr_wdata,_T_131}; // @[Cat.scala 30:58:@2939.8]
  assign _GEN_110 = _T_551 ? _T_1261 : _GEN_81; // @[rvcsr.scala 470:58:@2937.6]
  assign _T_1263 = {csr_wdata,_T_133}; // @[Cat.scala 30:58:@2944.8]
  assign _GEN_111 = _T_555 ? _T_1263 : _GEN_82; // @[rvcsr.scala 470:58:@2942.6]
  assign _T_1265 = {csr_wdata,_T_135}; // @[Cat.scala 30:58:@2949.8]
  assign _GEN_112 = _T_559 ? _T_1265 : _GEN_83; // @[rvcsr.scala 470:58:@2947.6]
  assign _T_1267 = {csr_wdata,_T_137}; // @[Cat.scala 30:58:@2954.8]
  assign _GEN_113 = _T_563 ? _T_1267 : _GEN_84; // @[rvcsr.scala 470:58:@2952.6]
  assign _T_1269 = {csr_wdata,_T_139}; // @[Cat.scala 30:58:@2959.8]
  assign _GEN_114 = _T_567 ? _T_1269 : _GEN_85; // @[rvcsr.scala 470:58:@2957.6]
  assign _T_1271 = {csr_wdata,_T_141}; // @[Cat.scala 30:58:@2964.8]
  assign _GEN_115 = _T_571 ? _T_1271 : _GEN_86; // @[rvcsr.scala 470:58:@2962.6]
  assign _T_1273 = {csr_wdata,_T_143}; // @[Cat.scala 30:58:@2969.8]
  assign _GEN_116 = _T_575 ? _T_1273 : _GEN_87; // @[rvcsr.scala 470:58:@2967.6]
  assign _T_1275 = {csr_wdata,_T_145}; // @[Cat.scala 30:58:@2974.8]
  assign _GEN_117 = _T_579 ? _T_1275 : _GEN_88; // @[rvcsr.scala 470:58:@2972.6]
  assign _T_1277 = {csr_wdata,_T_147}; // @[Cat.scala 30:58:@2979.8]
  assign _GEN_118 = _T_583 ? _T_1277 : _GEN_89; // @[rvcsr.scala 470:58:@2977.6]
  assign _T_1279 = {csr_wdata,_T_149}; // @[Cat.scala 30:58:@2984.8]
  assign _GEN_119 = _T_587 ? _T_1279 : _GEN_90; // @[rvcsr.scala 470:58:@2982.6]
  assign _T_1281 = {csr_wdata,_T_151}; // @[Cat.scala 30:58:@2989.8]
  assign _GEN_120 = _T_591 ? _T_1281 : _GEN_91; // @[rvcsr.scala 470:58:@2987.6]
  assign _T_1283 = {csr_wdata,_T_153}; // @[Cat.scala 30:58:@2994.8]
  assign _GEN_121 = _T_595 ? _T_1283 : _GEN_92; // @[rvcsr.scala 470:58:@2992.6]
  assign _T_1285 = {csr_wdata,_T_155}; // @[Cat.scala 30:58:@2999.8]
  assign _GEN_122 = _T_599 ? _T_1285 : _GEN_93; // @[rvcsr.scala 470:58:@2997.6]
  assign _T_1287 = {csr_wdata,_T_157}; // @[Cat.scala 30:58:@3004.8]
  assign _GEN_123 = _T_603 ? _T_1287 : _GEN_94; // @[rvcsr.scala 470:58:@3002.6]
  assign _T_1289 = {csr_wdata,_T_159}; // @[Cat.scala 30:58:@3009.8]
  assign _GEN_124 = _T_607 ? _T_1289 : _GEN_95; // @[rvcsr.scala 470:58:@3007.6]
  assign _T_1291 = {csr_wdata,_T_161}; // @[Cat.scala 30:58:@3014.8]
  assign _GEN_125 = _T_611 ? _T_1291 : _GEN_96; // @[rvcsr.scala 470:58:@3012.6]
  assign _T_1293 = {csr_wdata,_T_163}; // @[Cat.scala 30:58:@3019.8]
  assign _GEN_126 = _T_615 ? _T_1293 : _GEN_97; // @[rvcsr.scala 470:58:@3017.6]
  assign _T_1295 = {csr_wdata,_T_165}; // @[Cat.scala 30:58:@3024.8]
  assign _GEN_127 = _T_619 ? _T_1295 : _GEN_98; // @[rvcsr.scala 470:58:@3022.6]
  assign _T_1297 = {csr_wdata,_T_167}; // @[Cat.scala 30:58:@3029.8]
  assign _GEN_128 = _T_623 ? _T_1297 : _GEN_99; // @[rvcsr.scala 470:58:@3027.6]
  assign _T_1299 = {csr_wdata,_T_169}; // @[Cat.scala 30:58:@3034.8]
  assign _GEN_129 = _T_627 ? _T_1299 : _GEN_100; // @[rvcsr.scala 470:58:@3032.6]
  assign _T_1301 = {csr_wdata,_T_171}; // @[Cat.scala 30:58:@3039.8]
  assign _GEN_130 = _T_631 ? _T_1301 : _GEN_101; // @[rvcsr.scala 470:58:@3037.6]
  assign _GEN_131 = _T_633 ? csr_wdata : reg_mhpmevents_0; // @[rvcsr.scala 477:55:@3042.6]
  assign _GEN_132 = _T_635 ? csr_wdata : reg_mhpmevents_1; // @[rvcsr.scala 477:55:@3045.6]
  assign _GEN_133 = _T_637 ? csr_wdata : reg_mhpmevents_2; // @[rvcsr.scala 477:55:@3048.6]
  assign _GEN_134 = _T_639 ? csr_wdata : reg_mhpmevents_3; // @[rvcsr.scala 477:55:@3051.6]
  assign _GEN_135 = _T_641 ? csr_wdata : reg_mhpmevents_4; // @[rvcsr.scala 477:55:@3054.6]
  assign _GEN_136 = _T_643 ? csr_wdata : reg_mhpmevents_5; // @[rvcsr.scala 477:55:@3057.6]
  assign _GEN_137 = _T_645 ? csr_wdata : reg_mhpmevents_6; // @[rvcsr.scala 477:55:@3060.6]
  assign _GEN_138 = _T_647 ? csr_wdata : reg_mhpmevents_7; // @[rvcsr.scala 477:55:@3063.6]
  assign _GEN_139 = _T_649 ? csr_wdata : reg_mhpmevents_8; // @[rvcsr.scala 477:55:@3066.6]
  assign _GEN_140 = _T_651 ? csr_wdata : reg_mhpmevents_9; // @[rvcsr.scala 477:55:@3069.6]
  assign _GEN_141 = _T_653 ? csr_wdata : reg_mhpmevents_10; // @[rvcsr.scala 477:55:@3072.6]
  assign _GEN_142 = _T_655 ? csr_wdata : reg_mhpmevents_11; // @[rvcsr.scala 477:55:@3075.6]
  assign _GEN_143 = _T_657 ? csr_wdata : reg_mhpmevents_12; // @[rvcsr.scala 477:55:@3078.6]
  assign _GEN_144 = _T_659 ? csr_wdata : reg_mhpmevents_13; // @[rvcsr.scala 477:55:@3081.6]
  assign _GEN_145 = _T_661 ? csr_wdata : reg_mhpmevents_14; // @[rvcsr.scala 477:55:@3084.6]
  assign _GEN_146 = _T_663 ? csr_wdata : reg_mhpmevents_15; // @[rvcsr.scala 477:55:@3087.6]
  assign _GEN_147 = _T_665 ? csr_wdata : reg_mhpmevents_16; // @[rvcsr.scala 477:55:@3090.6]
  assign _GEN_148 = _T_667 ? csr_wdata : reg_mhpmevents_17; // @[rvcsr.scala 477:55:@3093.6]
  assign _GEN_149 = _T_669 ? csr_wdata : reg_mhpmevents_18; // @[rvcsr.scala 477:55:@3096.6]
  assign _GEN_150 = _T_671 ? csr_wdata : reg_mhpmevents_19; // @[rvcsr.scala 477:55:@3099.6]
  assign _GEN_151 = _T_673 ? csr_wdata : reg_mhpmevents_20; // @[rvcsr.scala 477:55:@3102.6]
  assign _GEN_152 = _T_675 ? csr_wdata : reg_mhpmevents_21; // @[rvcsr.scala 477:55:@3105.6]
  assign _GEN_153 = _T_677 ? csr_wdata : reg_mhpmevents_22; // @[rvcsr.scala 477:55:@3108.6]
  assign _GEN_154 = _T_679 ? csr_wdata : reg_mhpmevents_23; // @[rvcsr.scala 477:55:@3111.6]
  assign _GEN_155 = _T_681 ? csr_wdata : reg_mhpmevents_24; // @[rvcsr.scala 477:55:@3114.6]
  assign _GEN_156 = _T_683 ? csr_wdata : reg_mhpmevents_25; // @[rvcsr.scala 477:55:@3117.6]
  assign _GEN_157 = _T_685 ? csr_wdata : reg_mhpmevents_26; // @[rvcsr.scala 477:55:@3120.6]
  assign _GEN_158 = _T_687 ? csr_wdata : reg_mhpmevents_27; // @[rvcsr.scala 477:55:@3123.6]
  assign _GEN_159 = _T_689 ? csr_wdata : reg_mhpmevents_28; // @[rvcsr.scala 477:55:@3126.6]
  assign _T_1303 = {_T_113,csr_wdata}; // @[Cat.scala 30:58:@3131.8]
  assign _GEN_160 = _T_501 ? _T_1303 : _GEN_1; // @[rvcsr.scala 482:39:@3129.6]
  assign _T_1305 = {_T_112,csr_wdata}; // @[Cat.scala 30:58:@3136.8]
  assign _GEN_161 = _T_503 ? _T_1305 : reg_mtimecmp; // @[rvcsr.scala 487:42:@3134.6]
  assign _T_1307 = {csr_wdata,_T_111}; // @[Cat.scala 30:58:@3141.8]
  assign _GEN_162 = _T_505 ? _T_1307 : _GEN_160; // @[rvcsr.scala 492:40:@3139.6]
  assign _T_1308 = reg_mtimecmp[31:0]; // @[rvcsr.scala 499:56:@3145.8]
  assign _T_1309 = {csr_wdata,_T_1308}; // @[Cat.scala 30:58:@3146.8]
  assign _GEN_163 = _T_507 ? _T_1309 : _GEN_161; // @[rvcsr.scala 497:43:@3144.6]
  assign _GEN_164 = _T_473 ? csr_wdata : reg_medeleg; // @[rvcsr.scala 502:41:@3149.6]
  assign _GEN_165 = _T_475 ? csr_wdata : reg_mideleg; // @[rvcsr.scala 506:41:@3152.6]
  assign dcsr_rsrvd3 = reset ? 3'h0 : _T_385; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_166 = _T_509 ? _T_1065 : _T_384; // @[rvcsr.scala 510:38:@3155.6]
  assign _GEN_251 = csr_wen ? _GEN_166 : _T_384; // @[rvcsr.scala 393:19:@2545.4]
  assign dcsr_step = reset ? 1'h0 : _GEN_251; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_1328 = {dcsr_rsrvd3,dcsr_step}; // @[rvcsr.scala 514:30:@3187.8]
  assign _T_1329 = {_T_1328,dcsr_prv}; // @[rvcsr.scala 514:30:@3188.8]
  assign dcsr_stopcount = reset ? 1'h0 : _T_388; // @[rvcsr.scala 531:26:@3212.4]
  assign dcsr_stoptime = reset ? 1'h0 : _T_387; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_1330 = {dcsr_stopcount,dcsr_stoptime}; // @[rvcsr.scala 514:30:@3189.8]
  assign dcsr_cause = reset ? 3'h0 : _T_386; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_1331 = {_T_1330,dcsr_cause}; // @[rvcsr.scala 514:30:@3190.8]
  assign _T_1332 = {_T_1331,_T_1329}; // @[rvcsr.scala 514:30:@3191.8]
  assign dcsr_ebreaks = reset ? 1'h0 : _T_391; // @[rvcsr.scala 531:26:@3212.4]
  assign dcsr_ebreaku = reset ? 1'h0 : _T_390; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_1333 = {dcsr_ebreaks,dcsr_ebreaku}; // @[rvcsr.scala 514:30:@3192.8]
  assign dcsr_rsrvd2 = reset ? 1'h0 : _T_389; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_1334 = {_T_1333,dcsr_rsrvd2}; // @[rvcsr.scala 514:30:@3193.8]
  assign dcsr_ebreakh = reset ? 1'h0 : _T_392; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_1335 = {dcsr_ebreakm,dcsr_ebreakh}; // @[rvcsr.scala 514:30:@3194.8]
  assign dcsr_xdebugver = reset ? 4'h4 : _T_395; // @[rvcsr.scala 531:26:@3212.4]
  assign dcsr_rsrvd1 = reset ? 12'h0 : _T_394; // @[rvcsr.scala 531:26:@3212.4]
  assign _T_1336 = {dcsr_xdebugver,dcsr_rsrvd1}; // @[rvcsr.scala 514:30:@3195.8]
  assign _T_1337 = {_T_1336,_T_1335}; // @[rvcsr.scala 514:30:@3196.8]
  assign _T_1338 = {_T_1337,_T_1334}; // @[rvcsr.scala 514:30:@3197.8]
  assign _T_1339 = {_T_1338,_T_1332}; // @[rvcsr.scala 514:30:@3198.8]
  assign _GEN_168 = _T_509 ? _T_1339 : reg_dcsr; // @[rvcsr.scala 510:38:@3155.6]
  assign _GEN_169 = _T_511 ? csr_wdata : reg_dpc; // @[rvcsr.scala 517:37:@3201.6]
  assign _GEN_170 = _T_513 ? csr_wdata : reg_dscratch0; // @[rvcsr.scala 521:43:@3204.6]
  assign _GEN_171 = _T_515 ? csr_wdata : reg_dscratch1; // @[rvcsr.scala 525:43:@3207.6]
  assign _GEN_174 = csr_wen ? _GEN_56 : _GEN_38; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_177 = csr_wen ? _GEN_59 : reg_mie; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_178 = csr_wen ? _GEN_60 : reg_mtvec; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_179 = csr_wen ? _GEN_61 : reg_mcounteren; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_180 = csr_wen ? _GEN_62 : reg_mscratch; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_181 = csr_wen ? _GEN_63 : _GEN_52; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_182 = csr_wen ? _GEN_64 : _GEN_51; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_183 = csr_wen ? _GEN_65 : reg_mtval; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_186 = csr_wen ? _GEN_68 : _GEN_33; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_187 = csr_wen ? _GEN_71 : _GEN_0; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_188 = csr_wen ? _GEN_72 : _GEN_2; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_189 = csr_wen ? _GEN_102 : _GEN_3; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_190 = csr_wen ? _GEN_103 : _GEN_4; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_191 = csr_wen ? _GEN_104 : _GEN_5; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_192 = csr_wen ? _GEN_105 : _GEN_6; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_193 = csr_wen ? _GEN_106 : _GEN_7; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_194 = csr_wen ? _GEN_107 : _GEN_8; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_195 = csr_wen ? _GEN_108 : _GEN_9; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_196 = csr_wen ? _GEN_109 : _GEN_10; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_197 = csr_wen ? _GEN_110 : _GEN_11; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_198 = csr_wen ? _GEN_111 : _GEN_12; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_199 = csr_wen ? _GEN_112 : _GEN_13; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_200 = csr_wen ? _GEN_113 : _GEN_14; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_201 = csr_wen ? _GEN_114 : _GEN_15; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_202 = csr_wen ? _GEN_115 : _GEN_16; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_203 = csr_wen ? _GEN_116 : _GEN_17; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_204 = csr_wen ? _GEN_117 : _GEN_18; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_205 = csr_wen ? _GEN_118 : _GEN_19; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_206 = csr_wen ? _GEN_119 : _GEN_20; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_207 = csr_wen ? _GEN_120 : _GEN_21; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_208 = csr_wen ? _GEN_121 : _GEN_22; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_209 = csr_wen ? _GEN_122 : _GEN_23; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_210 = csr_wen ? _GEN_123 : _GEN_24; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_211 = csr_wen ? _GEN_124 : _GEN_25; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_212 = csr_wen ? _GEN_125 : _GEN_26; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_213 = csr_wen ? _GEN_126 : _GEN_27; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_214 = csr_wen ? _GEN_127 : _GEN_28; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_215 = csr_wen ? _GEN_128 : _GEN_29; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_216 = csr_wen ? _GEN_129 : _GEN_30; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_217 = csr_wen ? _GEN_130 : _GEN_31; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_218 = csr_wen ? _GEN_131 : reg_mhpmevents_0; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_219 = csr_wen ? _GEN_132 : reg_mhpmevents_1; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_220 = csr_wen ? _GEN_133 : reg_mhpmevents_2; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_221 = csr_wen ? _GEN_134 : reg_mhpmevents_3; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_222 = csr_wen ? _GEN_135 : reg_mhpmevents_4; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_223 = csr_wen ? _GEN_136 : reg_mhpmevents_5; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_224 = csr_wen ? _GEN_137 : reg_mhpmevents_6; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_225 = csr_wen ? _GEN_138 : reg_mhpmevents_7; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_226 = csr_wen ? _GEN_139 : reg_mhpmevents_8; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_227 = csr_wen ? _GEN_140 : reg_mhpmevents_9; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_228 = csr_wen ? _GEN_141 : reg_mhpmevents_10; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_229 = csr_wen ? _GEN_142 : reg_mhpmevents_11; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_230 = csr_wen ? _GEN_143 : reg_mhpmevents_12; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_231 = csr_wen ? _GEN_144 : reg_mhpmevents_13; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_232 = csr_wen ? _GEN_145 : reg_mhpmevents_14; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_233 = csr_wen ? _GEN_146 : reg_mhpmevents_15; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_234 = csr_wen ? _GEN_147 : reg_mhpmevents_16; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_235 = csr_wen ? _GEN_148 : reg_mhpmevents_17; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_236 = csr_wen ? _GEN_149 : reg_mhpmevents_18; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_237 = csr_wen ? _GEN_150 : reg_mhpmevents_19; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_238 = csr_wen ? _GEN_151 : reg_mhpmevents_20; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_239 = csr_wen ? _GEN_152 : reg_mhpmevents_21; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_240 = csr_wen ? _GEN_153 : reg_mhpmevents_22; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_241 = csr_wen ? _GEN_154 : reg_mhpmevents_23; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_242 = csr_wen ? _GEN_155 : reg_mhpmevents_24; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_243 = csr_wen ? _GEN_156 : reg_mhpmevents_25; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_244 = csr_wen ? _GEN_157 : reg_mhpmevents_26; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_245 = csr_wen ? _GEN_158 : reg_mhpmevents_27; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_246 = csr_wen ? _GEN_159 : reg_mhpmevents_28; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_247 = csr_wen ? _GEN_162 : _GEN_1; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_248 = csr_wen ? _GEN_163 : reg_mtimecmp; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_249 = csr_wen ? _GEN_164 : reg_medeleg; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_250 = csr_wen ? _GEN_165 : reg_mideleg; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_253 = csr_wen ? _GEN_168 : reg_dcsr; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_254 = csr_wen ? _GEN_169 : reg_dpc; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_255 = csr_wen ? _GEN_170 : reg_dscratch0; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_256 = csr_wen ? _GEN_171 : reg_dscratch1; // @[rvcsr.scala 393:19:@2545.4]
  assign _GEN_257 = reset ? 2'h3 : _GEN_46; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_279 = reset ? _T_447 : _GEN_174; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_280 = reset ? 32'h100 : _GEN_178; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_281 = reset ? 32'h0 : _GEN_249; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_282 = reset ? 32'h0 : _GEN_250; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_283 = reset ? 32'h0 : _GEN_186; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_284 = reset ? 32'h0 : _GEN_177; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_285 = reset ? 64'h0 : _GEN_247; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_286 = reset ? 64'h0 : _GEN_248; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_287 = reset ? 64'h0 : _GEN_187; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_288 = reset ? 64'h0 : _GEN_188; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_289 = reset ? 64'h0 : _GEN_189; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_290 = reset ? 64'h0 : _GEN_190; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_291 = reset ? 64'h0 : _GEN_191; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_292 = reset ? 64'h0 : _GEN_192; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_293 = reset ? 64'h0 : _GEN_193; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_294 = reset ? 64'h0 : _GEN_194; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_295 = reset ? 64'h0 : _GEN_195; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_296 = reset ? 64'h0 : _GEN_196; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_297 = reset ? 64'h0 : _GEN_197; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_298 = reset ? 64'h0 : _GEN_198; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_299 = reset ? 64'h0 : _GEN_199; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_300 = reset ? 64'h0 : _GEN_200; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_301 = reset ? 64'h0 : _GEN_201; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_302 = reset ? 64'h0 : _GEN_202; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_303 = reset ? 64'h0 : _GEN_203; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_304 = reset ? 64'h0 : _GEN_204; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_305 = reset ? 64'h0 : _GEN_205; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_306 = reset ? 64'h0 : _GEN_206; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_307 = reset ? 64'h0 : _GEN_207; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_308 = reset ? 64'h0 : _GEN_208; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_309 = reset ? 64'h0 : _GEN_209; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_310 = reset ? 64'h0 : _GEN_210; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_311 = reset ? 64'h0 : _GEN_211; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_312 = reset ? 64'h0 : _GEN_212; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_313 = reset ? 64'h0 : _GEN_213; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_314 = reset ? 64'h0 : _GEN_214; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_315 = reset ? 64'h0 : _GEN_215; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_316 = reset ? 64'h0 : _GEN_216; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_317 = reset ? 64'h0 : _GEN_217; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_318 = reset ? 32'h0 : _GEN_218; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_319 = reset ? 32'h0 : _GEN_219; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_320 = reset ? 32'h0 : _GEN_220; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_321 = reset ? 32'h0 : _GEN_221; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_322 = reset ? 32'h0 : _GEN_222; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_323 = reset ? 32'h0 : _GEN_223; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_324 = reset ? 32'h0 : _GEN_224; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_325 = reset ? 32'h0 : _GEN_225; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_326 = reset ? 32'h0 : _GEN_226; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_327 = reset ? 32'h0 : _GEN_227; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_328 = reset ? 32'h0 : _GEN_228; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_329 = reset ? 32'h0 : _GEN_229; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_330 = reset ? 32'h0 : _GEN_230; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_331 = reset ? 32'h0 : _GEN_231; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_332 = reset ? 32'h0 : _GEN_232; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_333 = reset ? 32'h0 : _GEN_233; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_334 = reset ? 32'h0 : _GEN_234; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_335 = reset ? 32'h0 : _GEN_235; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_336 = reset ? 32'h0 : _GEN_236; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_337 = reset ? 32'h0 : _GEN_237; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_338 = reset ? 32'h0 : _GEN_238; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_339 = reset ? 32'h0 : _GEN_239; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_340 = reset ? 32'h0 : _GEN_240; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_341 = reset ? 32'h0 : _GEN_241; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_342 = reset ? 32'h0 : _GEN_242; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_343 = reset ? 32'h0 : _GEN_243; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_344 = reset ? 32'h0 : _GEN_244; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_345 = reset ? 32'h0 : _GEN_245; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_346 = reset ? 32'h0 : _GEN_246; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_347 = reset ? 32'h0 : _GEN_179; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_348 = reset ? 32'h0 : _GEN_180; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_349 = reset ? 32'h0 : _GEN_181; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_350 = reset ? 32'h0 : _GEN_182; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_351 = reset ? 32'h0 : _GEN_183; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_366 = reset ? _T_1339 : _GEN_253; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_367 = reset ? 32'h0 : _GEN_254; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_368 = reset ? 32'h0 : _GEN_255; // @[rvcsr.scala 531:26:@3212.4]
  assign _GEN_369 = reset ? 32'h0 : _GEN_256; // @[rvcsr.scala 531:26:@3212.4]
  assign io_rdata = _T_1044;
  assign io_csr_excp = _T_406;
  assign io_csr_evec = _GEN_53;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  reg_priv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  reg_mstatus = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  reg_mtvec = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  reg_medeleg = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  reg_mideleg = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  reg_mip = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  reg_mie = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{$random}};
  reg_mtime = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{$random}};
  reg_mtimecmp = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{$random}};
  reg_mcycle = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{$random}};
  reg_minstret = _RAND_10[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{$random}};
  reg_mhpmcounters_0 = _RAND_11[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{$random}};
  reg_mhpmcounters_1 = _RAND_12[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{$random}};
  reg_mhpmcounters_2 = _RAND_13[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{$random}};
  reg_mhpmcounters_3 = _RAND_14[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{$random}};
  reg_mhpmcounters_4 = _RAND_15[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{$random}};
  reg_mhpmcounters_5 = _RAND_16[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{$random}};
  reg_mhpmcounters_6 = _RAND_17[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{$random}};
  reg_mhpmcounters_7 = _RAND_18[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{$random}};
  reg_mhpmcounters_8 = _RAND_19[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{$random}};
  reg_mhpmcounters_9 = _RAND_20[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{$random}};
  reg_mhpmcounters_10 = _RAND_21[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{$random}};
  reg_mhpmcounters_11 = _RAND_22[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{$random}};
  reg_mhpmcounters_12 = _RAND_23[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{$random}};
  reg_mhpmcounters_13 = _RAND_24[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{$random}};
  reg_mhpmcounters_14 = _RAND_25[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{$random}};
  reg_mhpmcounters_15 = _RAND_26[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{$random}};
  reg_mhpmcounters_16 = _RAND_27[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{$random}};
  reg_mhpmcounters_17 = _RAND_28[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{$random}};
  reg_mhpmcounters_18 = _RAND_29[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{$random}};
  reg_mhpmcounters_19 = _RAND_30[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{$random}};
  reg_mhpmcounters_20 = _RAND_31[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{$random}};
  reg_mhpmcounters_21 = _RAND_32[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{$random}};
  reg_mhpmcounters_22 = _RAND_33[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{$random}};
  reg_mhpmcounters_23 = _RAND_34[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{$random}};
  reg_mhpmcounters_24 = _RAND_35[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{$random}};
  reg_mhpmcounters_25 = _RAND_36[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{$random}};
  reg_mhpmcounters_26 = _RAND_37[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{$random}};
  reg_mhpmcounters_27 = _RAND_38[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{$random}};
  reg_mhpmcounters_28 = _RAND_39[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  reg_mhpmevents_0 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  reg_mhpmevents_1 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  reg_mhpmevents_2 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  reg_mhpmevents_3 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  reg_mhpmevents_4 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  reg_mhpmevents_5 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  reg_mhpmevents_6 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  reg_mhpmevents_7 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  reg_mhpmevents_8 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  reg_mhpmevents_9 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  reg_mhpmevents_10 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  reg_mhpmevents_11 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  reg_mhpmevents_12 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  reg_mhpmevents_13 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  reg_mhpmevents_14 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  reg_mhpmevents_15 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  reg_mhpmevents_16 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  reg_mhpmevents_17 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  reg_mhpmevents_18 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  reg_mhpmevents_19 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  reg_mhpmevents_20 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  reg_mhpmevents_21 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  reg_mhpmevents_22 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  reg_mhpmevents_23 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  reg_mhpmevents_24 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  reg_mhpmevents_25 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  reg_mhpmevents_26 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  reg_mhpmevents_27 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  reg_mhpmevents_28 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  reg_mcounteren = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  reg_mscratch = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  reg_mepc = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  reg_mcause = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  reg_mtval = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  reg_dcsr = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  reg_dpc = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  reg_dscratch0 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  reg_dscratch1 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_priv <= 2'h3;
    end else begin
      if (_T_456) begin
        if (reset) begin
          reg_priv <= 2'h3;
        end else begin
          reg_priv <= _T_383;
        end
      end else begin
        if (_T_426) begin
          if (reset) begin
            reg_priv <= 2'h3;
          end else begin
            reg_priv <= _T_328;
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus <= _T_447;
    end else begin
      if (csr_wen) begin
        if (_T_469) begin
          reg_mstatus <= _T_447;
        end else begin
          if (_T_426) begin
            reg_mstatus <= _T_447;
          end
        end
      end else begin
        if (_T_426) begin
          reg_mstatus <= _T_447;
        end
      end
    end
    if (reset) begin
      reg_mtvec <= 32'h100;
    end else begin
      if (csr_wen) begin
        if (_T_479) begin
          reg_mtvec <= _T_1140;
        end
      end
    end
    if (reset) begin
      reg_medeleg <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_473) begin
          reg_medeleg <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mideleg <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_475) begin
          reg_mideleg <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mip <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_491) begin
          reg_mip <= {{1'd0}, _T_420};
        end else begin
          if (_T_407) begin
            reg_mip <= {{1'd0}, _T_420};
          end
        end
      end else begin
        if (_T_407) begin
          reg_mip <= {{1'd0}, _T_420};
        end
      end
    end
    if (reset) begin
      reg_mie <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_477) begin
          reg_mie <= {{1'd0}, _T_1133};
        end
      end
    end
    if (reset) begin
      reg_mtime <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_505) begin
          reg_mtime <= _T_1307;
        end else begin
          if (_T_501) begin
            reg_mtime <= _T_1303;
          end else begin
            if (counteren_TM) begin
              reg_mtime <= _T_220;
            end
          end
        end
      end else begin
        if (counteren_TM) begin
          reg_mtime <= _T_220;
        end
      end
    end
    if (reset) begin
      reg_mtimecmp <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_507) begin
          reg_mtimecmp <= _T_1309;
        end else begin
          if (_T_503) begin
            reg_mtimecmp <= _T_1305;
          end
        end
      end
    end
    if (reset) begin
      reg_mcycle <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_497) begin
          reg_mcycle <= _T_1183;
        end else begin
          if (_T_493) begin
            reg_mcycle <= _T_1179;
          end else begin
            if (counteren_CY) begin
              reg_mcycle <= _T_217;
            end
          end
        end
      end else begin
        if (counteren_CY) begin
          reg_mcycle <= _T_217;
        end
      end
    end
    if (reset) begin
      reg_minstret <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_499) begin
          reg_minstret <= _T_1185;
        end else begin
          if (_T_495) begin
            reg_minstret <= _T_1181;
          end else begin
            if (counteren_IR) begin
              reg_minstret <= _T_223;
            end
          end
        end
      end else begin
        if (counteren_IR) begin
          reg_minstret <= _T_223;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_0 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_519) begin
          reg_mhpmcounters_0 <= _T_1245;
        end else begin
          if (_T_517) begin
            reg_mhpmcounters_0 <= _T_1187;
          end else begin
            if (counteren_HPM_0) begin
              reg_mhpmcounters_0 <= _T_226;
            end
          end
        end
      end else begin
        if (counteren_HPM_0) begin
          reg_mhpmcounters_0 <= _T_226;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_1 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_523) begin
          reg_mhpmcounters_1 <= _T_1247;
        end else begin
          if (_T_521) begin
            reg_mhpmcounters_1 <= _T_1189;
          end else begin
            if (counteren_HPM_1) begin
              reg_mhpmcounters_1 <= _T_229;
            end
          end
        end
      end else begin
        if (counteren_HPM_1) begin
          reg_mhpmcounters_1 <= _T_229;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_2 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_527) begin
          reg_mhpmcounters_2 <= _T_1249;
        end else begin
          if (_T_525) begin
            reg_mhpmcounters_2 <= _T_1191;
          end else begin
            if (counteren_HPM_2) begin
              reg_mhpmcounters_2 <= _T_232;
            end
          end
        end
      end else begin
        if (counteren_HPM_2) begin
          reg_mhpmcounters_2 <= _T_232;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_3 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_531) begin
          reg_mhpmcounters_3 <= _T_1251;
        end else begin
          if (_T_529) begin
            reg_mhpmcounters_3 <= _T_1193;
          end else begin
            if (counteren_HPM_3) begin
              reg_mhpmcounters_3 <= _T_235;
            end
          end
        end
      end else begin
        if (counteren_HPM_3) begin
          reg_mhpmcounters_3 <= _T_235;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_4 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_535) begin
          reg_mhpmcounters_4 <= _T_1253;
        end else begin
          if (_T_533) begin
            reg_mhpmcounters_4 <= _T_1195;
          end else begin
            if (counteren_HPM_4) begin
              reg_mhpmcounters_4 <= _T_238;
            end
          end
        end
      end else begin
        if (counteren_HPM_4) begin
          reg_mhpmcounters_4 <= _T_238;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_5 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_539) begin
          reg_mhpmcounters_5 <= _T_1255;
        end else begin
          if (_T_537) begin
            reg_mhpmcounters_5 <= _T_1197;
          end else begin
            if (counteren_HPM_5) begin
              reg_mhpmcounters_5 <= _T_241;
            end
          end
        end
      end else begin
        if (counteren_HPM_5) begin
          reg_mhpmcounters_5 <= _T_241;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_6 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_543) begin
          reg_mhpmcounters_6 <= _T_1257;
        end else begin
          if (_T_541) begin
            reg_mhpmcounters_6 <= _T_1199;
          end else begin
            if (counteren_HPM_6) begin
              reg_mhpmcounters_6 <= _T_244;
            end
          end
        end
      end else begin
        if (counteren_HPM_6) begin
          reg_mhpmcounters_6 <= _T_244;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_7 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_547) begin
          reg_mhpmcounters_7 <= _T_1259;
        end else begin
          if (_T_545) begin
            reg_mhpmcounters_7 <= _T_1201;
          end else begin
            if (counteren_HPM_7) begin
              reg_mhpmcounters_7 <= _T_247;
            end
          end
        end
      end else begin
        if (counteren_HPM_7) begin
          reg_mhpmcounters_7 <= _T_247;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_8 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_551) begin
          reg_mhpmcounters_8 <= _T_1261;
        end else begin
          if (_T_549) begin
            reg_mhpmcounters_8 <= _T_1203;
          end else begin
            if (counteren_HPM_8) begin
              reg_mhpmcounters_8 <= _T_250;
            end
          end
        end
      end else begin
        if (counteren_HPM_8) begin
          reg_mhpmcounters_8 <= _T_250;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_9 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_555) begin
          reg_mhpmcounters_9 <= _T_1263;
        end else begin
          if (_T_553) begin
            reg_mhpmcounters_9 <= _T_1205;
          end else begin
            if (counteren_HPM_9) begin
              reg_mhpmcounters_9 <= _T_253;
            end
          end
        end
      end else begin
        if (counteren_HPM_9) begin
          reg_mhpmcounters_9 <= _T_253;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_10 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_559) begin
          reg_mhpmcounters_10 <= _T_1265;
        end else begin
          if (_T_557) begin
            reg_mhpmcounters_10 <= _T_1207;
          end else begin
            if (counteren_HPM_10) begin
              reg_mhpmcounters_10 <= _T_256;
            end
          end
        end
      end else begin
        if (counteren_HPM_10) begin
          reg_mhpmcounters_10 <= _T_256;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_11 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_563) begin
          reg_mhpmcounters_11 <= _T_1267;
        end else begin
          if (_T_561) begin
            reg_mhpmcounters_11 <= _T_1209;
          end else begin
            if (counteren_HPM_11) begin
              reg_mhpmcounters_11 <= _T_259;
            end
          end
        end
      end else begin
        if (counteren_HPM_11) begin
          reg_mhpmcounters_11 <= _T_259;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_12 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_567) begin
          reg_mhpmcounters_12 <= _T_1269;
        end else begin
          if (_T_565) begin
            reg_mhpmcounters_12 <= _T_1211;
          end else begin
            if (counteren_HPM_12) begin
              reg_mhpmcounters_12 <= _T_262;
            end
          end
        end
      end else begin
        if (counteren_HPM_12) begin
          reg_mhpmcounters_12 <= _T_262;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_13 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_571) begin
          reg_mhpmcounters_13 <= _T_1271;
        end else begin
          if (_T_569) begin
            reg_mhpmcounters_13 <= _T_1213;
          end else begin
            if (counteren_HPM_13) begin
              reg_mhpmcounters_13 <= _T_265;
            end
          end
        end
      end else begin
        if (counteren_HPM_13) begin
          reg_mhpmcounters_13 <= _T_265;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_14 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_575) begin
          reg_mhpmcounters_14 <= _T_1273;
        end else begin
          if (_T_573) begin
            reg_mhpmcounters_14 <= _T_1215;
          end else begin
            if (counteren_HPM_14) begin
              reg_mhpmcounters_14 <= _T_268;
            end
          end
        end
      end else begin
        if (counteren_HPM_14) begin
          reg_mhpmcounters_14 <= _T_268;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_15 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_579) begin
          reg_mhpmcounters_15 <= _T_1275;
        end else begin
          if (_T_577) begin
            reg_mhpmcounters_15 <= _T_1217;
          end else begin
            if (counteren_HPM_15) begin
              reg_mhpmcounters_15 <= _T_271;
            end
          end
        end
      end else begin
        if (counteren_HPM_15) begin
          reg_mhpmcounters_15 <= _T_271;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_16 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_583) begin
          reg_mhpmcounters_16 <= _T_1277;
        end else begin
          if (_T_581) begin
            reg_mhpmcounters_16 <= _T_1219;
          end else begin
            if (counteren_HPM_16) begin
              reg_mhpmcounters_16 <= _T_274;
            end
          end
        end
      end else begin
        if (counteren_HPM_16) begin
          reg_mhpmcounters_16 <= _T_274;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_17 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_587) begin
          reg_mhpmcounters_17 <= _T_1279;
        end else begin
          if (_T_585) begin
            reg_mhpmcounters_17 <= _T_1221;
          end else begin
            if (counteren_HPM_17) begin
              reg_mhpmcounters_17 <= _T_277;
            end
          end
        end
      end else begin
        if (counteren_HPM_17) begin
          reg_mhpmcounters_17 <= _T_277;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_18 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_591) begin
          reg_mhpmcounters_18 <= _T_1281;
        end else begin
          if (_T_589) begin
            reg_mhpmcounters_18 <= _T_1223;
          end else begin
            if (counteren_HPM_18) begin
              reg_mhpmcounters_18 <= _T_280;
            end
          end
        end
      end else begin
        if (counteren_HPM_18) begin
          reg_mhpmcounters_18 <= _T_280;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_19 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_595) begin
          reg_mhpmcounters_19 <= _T_1283;
        end else begin
          if (_T_593) begin
            reg_mhpmcounters_19 <= _T_1225;
          end else begin
            if (counteren_HPM_19) begin
              reg_mhpmcounters_19 <= _T_283;
            end
          end
        end
      end else begin
        if (counteren_HPM_19) begin
          reg_mhpmcounters_19 <= _T_283;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_20 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_599) begin
          reg_mhpmcounters_20 <= _T_1285;
        end else begin
          if (_T_597) begin
            reg_mhpmcounters_20 <= _T_1227;
          end else begin
            if (counteren_HPM_20) begin
              reg_mhpmcounters_20 <= _T_286;
            end
          end
        end
      end else begin
        if (counteren_HPM_20) begin
          reg_mhpmcounters_20 <= _T_286;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_21 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_603) begin
          reg_mhpmcounters_21 <= _T_1287;
        end else begin
          if (_T_601) begin
            reg_mhpmcounters_21 <= _T_1229;
          end else begin
            if (counteren_HPM_21) begin
              reg_mhpmcounters_21 <= _T_289;
            end
          end
        end
      end else begin
        if (counteren_HPM_21) begin
          reg_mhpmcounters_21 <= _T_289;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_22 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_607) begin
          reg_mhpmcounters_22 <= _T_1289;
        end else begin
          if (_T_605) begin
            reg_mhpmcounters_22 <= _T_1231;
          end else begin
            if (counteren_HPM_22) begin
              reg_mhpmcounters_22 <= _T_292;
            end
          end
        end
      end else begin
        if (counteren_HPM_22) begin
          reg_mhpmcounters_22 <= _T_292;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_23 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_611) begin
          reg_mhpmcounters_23 <= _T_1291;
        end else begin
          if (_T_609) begin
            reg_mhpmcounters_23 <= _T_1233;
          end else begin
            if (counteren_HPM_23) begin
              reg_mhpmcounters_23 <= _T_295;
            end
          end
        end
      end else begin
        if (counteren_HPM_23) begin
          reg_mhpmcounters_23 <= _T_295;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_24 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_615) begin
          reg_mhpmcounters_24 <= _T_1293;
        end else begin
          if (_T_613) begin
            reg_mhpmcounters_24 <= _T_1235;
          end else begin
            if (counteren_HPM_24) begin
              reg_mhpmcounters_24 <= _T_298;
            end
          end
        end
      end else begin
        if (counteren_HPM_24) begin
          reg_mhpmcounters_24 <= _T_298;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_25 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_619) begin
          reg_mhpmcounters_25 <= _T_1295;
        end else begin
          if (_T_617) begin
            reg_mhpmcounters_25 <= _T_1237;
          end else begin
            if (counteren_HPM_25) begin
              reg_mhpmcounters_25 <= _T_301;
            end
          end
        end
      end else begin
        if (counteren_HPM_25) begin
          reg_mhpmcounters_25 <= _T_301;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_26 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_623) begin
          reg_mhpmcounters_26 <= _T_1297;
        end else begin
          if (_T_621) begin
            reg_mhpmcounters_26 <= _T_1239;
          end else begin
            if (counteren_HPM_26) begin
              reg_mhpmcounters_26 <= _T_304;
            end
          end
        end
      end else begin
        if (counteren_HPM_26) begin
          reg_mhpmcounters_26 <= _T_304;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_27 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_627) begin
          reg_mhpmcounters_27 <= _T_1299;
        end else begin
          if (_T_625) begin
            reg_mhpmcounters_27 <= _T_1241;
          end else begin
            if (counteren_HPM_27) begin
              reg_mhpmcounters_27 <= _T_307;
            end
          end
        end
      end else begin
        if (counteren_HPM_27) begin
          reg_mhpmcounters_27 <= _T_307;
        end
      end
    end
    if (reset) begin
      reg_mhpmcounters_28 <= 64'h0;
    end else begin
      if (csr_wen) begin
        if (_T_631) begin
          reg_mhpmcounters_28 <= _T_1301;
        end else begin
          if (_T_629) begin
            reg_mhpmcounters_28 <= _T_1243;
          end else begin
            if (counteren_HPM_28) begin
              reg_mhpmcounters_28 <= _T_310;
            end
          end
        end
      end else begin
        if (counteren_HPM_28) begin
          reg_mhpmcounters_28 <= _T_310;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_0 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_633) begin
          reg_mhpmevents_0 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_1 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_635) begin
          reg_mhpmevents_1 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_2 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_637) begin
          reg_mhpmevents_2 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_3 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_639) begin
          reg_mhpmevents_3 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_4 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_641) begin
          reg_mhpmevents_4 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_5 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_643) begin
          reg_mhpmevents_5 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_6 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_645) begin
          reg_mhpmevents_6 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_7 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_647) begin
          reg_mhpmevents_7 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_8 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_649) begin
          reg_mhpmevents_8 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_9 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_651) begin
          reg_mhpmevents_9 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_10 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_653) begin
          reg_mhpmevents_10 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_11 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_655) begin
          reg_mhpmevents_11 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_12 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_657) begin
          reg_mhpmevents_12 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_13 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_659) begin
          reg_mhpmevents_13 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_14 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_661) begin
          reg_mhpmevents_14 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_15 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_663) begin
          reg_mhpmevents_15 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_16 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_665) begin
          reg_mhpmevents_16 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_17 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_667) begin
          reg_mhpmevents_17 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_18 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_669) begin
          reg_mhpmevents_18 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_19 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_671) begin
          reg_mhpmevents_19 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_20 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_673) begin
          reg_mhpmevents_20 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_21 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_675) begin
          reg_mhpmevents_21 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_22 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_677) begin
          reg_mhpmevents_22 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_23 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_679) begin
          reg_mhpmevents_23 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_24 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_681) begin
          reg_mhpmevents_24 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_25 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_683) begin
          reg_mhpmevents_25 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_26 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_685) begin
          reg_mhpmevents_26 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_27 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_687) begin
          reg_mhpmevents_27 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mhpmevents_28 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_689) begin
          reg_mhpmevents_28 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mcounteren <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_481) begin
          reg_mcounteren <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mscratch <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_483) begin
          reg_mscratch <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_mepc <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_485) begin
          reg_mepc <= _T_1140;
        end else begin
          if (io_core_excp) begin
            if (_T_458) begin
              reg_mepc <= io_core_pc;
            end
          end
        end
      end else begin
        if (io_core_excp) begin
          if (_T_458) begin
            reg_mepc <= io_core_pc;
          end
        end
      end
    end
    if (reset) begin
      reg_mcause <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_487) begin
          reg_mcause <= csr_wdata;
        end else begin
          if (io_core_excp) begin
            if (_T_458) begin
              reg_mcause <= {{28'd0}, io_core_cause};
            end else begin
              if (inst_ebreak) begin
                reg_mcause <= 32'h3;
              end else begin
                if (inst_ecall) begin
                  reg_mcause <= 32'hb;
                end
              end
            end
          end else begin
            if (inst_ebreak) begin
              reg_mcause <= 32'h3;
            end else begin
              if (inst_ecall) begin
                reg_mcause <= 32'hb;
              end
            end
          end
        end
      end else begin
        if (io_core_excp) begin
          if (_T_458) begin
            reg_mcause <= {{28'd0}, io_core_cause};
          end else begin
            if (inst_ebreak) begin
              reg_mcause <= 32'h3;
            end else begin
              if (inst_ecall) begin
                reg_mcause <= 32'hb;
              end
            end
          end
        end else begin
          if (inst_ebreak) begin
            reg_mcause <= 32'h3;
          end else begin
            if (inst_ecall) begin
              reg_mcause <= 32'hb;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mtval <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_489) begin
          reg_mtval <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_dcsr <= _T_1339;
    end else begin
      if (csr_wen) begin
        if (_T_509) begin
          reg_dcsr <= _T_1339;
        end
      end
    end
    if (reset) begin
      reg_dpc <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_511) begin
          reg_dpc <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_dscratch0 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_513) begin
          reg_dscratch0 <= csr_wdata;
        end
      end
    end
    if (reset) begin
      reg_dscratch1 <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_515) begin
          reg_dscratch1 <= csr_wdata;
        end
      end
    end
  end
endmodule
module rvdpath( // @[:@3439.2]
  input         clock, // @[:@3440.4]
  input         reset, // @[:@3441.4]
  output [31:0] io_imem_req_addr, // @[:@3442.4]
  output        io_imem_req_valid, // @[:@3442.4]
  input  [31:0] io_imem_resp_data, // @[:@3442.4]
  input         io_imem_resp_valid, // @[:@3442.4]
  output [31:0] io_dmem_req_addr, // @[:@3442.4]
  output [31:0] io_dmem_req_data, // @[:@3442.4]
  output        io_dmem_req_mfunc, // @[:@3442.4]
  output [1:0]  io_dmem_req_mtype, // @[:@3442.4]
  output        io_dmem_req_valid, // @[:@3442.4]
  input         io_dmem_req_ready, // @[:@3442.4]
  input  [31:0] io_dmem_resp_data, // @[:@3442.4]
  input         io_dmem_resp_valid, // @[:@3442.4]
  output [31:0] io_d2c_inst, // @[:@3442.4]
  output        io_d2c_dexcp, // @[:@3442.4]
  input  [3:0]  io_c2d_alu_func, // @[:@3442.4]
  input  [2:0]  io_c2d_op2_sel, // @[:@3442.4]
  input         io_c2d_reg_wren, // @[:@3442.4]
  input         io_c2d_mem_wren, // @[:@3442.4]
  input         io_c2d_mem_en, // @[:@3442.4]
  input  [1:0]  io_c2d_wb_sel, // @[:@3442.4]
  input  [2:0]  io_c2d_mem_type, // @[:@3442.4]
  input  [1:0]  io_c2d_pc_sel, // @[:@3442.4]
  input  [2:0]  io_c2d_br_sel, // @[:@3442.4]
  input  [1:0]  io_c2d_op1_sel, // @[:@3442.4]
  input  [2:0]  io_c2d_csr_cmd, // @[:@3442.4]
  input         io_c2d_cexcp, // @[:@3442.4]
  input  [3:0]  io_c2d_ccause, // @[:@3442.4]
  input  [4:0]  io_ddpath_addr, // @[:@3442.4]
  input  [31:0] io_ddpath_wdata, // @[:@3442.4]
  input         io_ddpath_valid, // @[:@3442.4]
  output [31:0] io_ddpath_rdata // @[:@3442.4]
);
  reg [31:0] pc; // @[rvdpath.scala 44:17:@3480.4]
  reg [31:0] _RAND_0;
  reg [31:0] regfile_0; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_1;
  reg [31:0] regfile_1; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_2;
  reg [31:0] regfile_2; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_3;
  reg [31:0] regfile_3; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_4;
  reg [31:0] regfile_4; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_5;
  reg [31:0] regfile_5; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_6;
  reg [31:0] regfile_6; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_7;
  reg [31:0] regfile_7; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_8;
  reg [31:0] regfile_8; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_9;
  reg [31:0] regfile_9; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_10;
  reg [31:0] regfile_10; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_11;
  reg [31:0] regfile_11; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_12;
  reg [31:0] regfile_12; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_13;
  reg [31:0] regfile_13; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_14;
  reg [31:0] regfile_14; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_15;
  reg [31:0] regfile_15; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_16;
  reg [31:0] regfile_16; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_17;
  reg [31:0] regfile_17; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_18;
  reg [31:0] regfile_18; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_19;
  reg [31:0] regfile_19; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_20;
  reg [31:0] regfile_20; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_21;
  reg [31:0] regfile_21; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_22;
  reg [31:0] regfile_22; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_23;
  reg [31:0] regfile_23; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_24;
  reg [31:0] regfile_24; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_25;
  reg [31:0] regfile_25; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_26;
  reg [31:0] regfile_26; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_27;
  reg [31:0] regfile_27; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_28;
  reg [31:0] regfile_28; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_29;
  reg [31:0] regfile_29; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_30;
  reg [31:0] regfile_30; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_31;
  reg [31:0] regfile_31; // @[rvdpath.scala 96:22:@3518.4]
  reg [31:0] _RAND_32;
  wire  csr_clock; // @[rvdpath.scala 251:21:@3741.4]
  wire  csr_reset; // @[rvdpath.scala 251:21:@3741.4]
  wire [11:0] csr_io_addr; // @[rvdpath.scala 251:21:@3741.4]
  wire [31:0] csr_io_wdata; // @[rvdpath.scala 251:21:@3741.4]
  wire [31:0] csr_io_rdata; // @[rvdpath.scala 251:21:@3741.4]
  wire [2:0] csr_io_op; // @[rvdpath.scala 251:21:@3741.4]
  wire [31:0] csr_io_core_pc; // @[rvdpath.scala 251:21:@3741.4]
  wire  csr_io_core_excp; // @[rvdpath.scala 251:21:@3741.4]
  wire [3:0] csr_io_core_cause; // @[rvdpath.scala 251:21:@3741.4]
  wire  csr_io_csr_excp; // @[rvdpath.scala 251:21:@3741.4]
  wire [31:0] csr_io_csr_evec; // @[rvdpath.scala 251:21:@3741.4]
  wire [32:0] _T_71; // @[rvdpath.scala 52:17:@3486.4]
  wire [31:0] pc_a4; // @[rvdpath.scala 52:17:@3487.4]
  wire  _T_73; // @[Mux.scala 46:19:@3489.4]
  wire [31:0] pc_ex; // @[rvdpath.scala 50:21:@3485.4]
  wire [31:0] _T_74; // @[Mux.scala 46:16:@3490.4]
  wire  _T_75; // @[Mux.scala 46:19:@3491.4]
  wire  _T_261; // @[Mux.scala 46:19:@3638.4]
  wire  _T_197; // @[Mux.scala 46:19:@3571.4]
  wire [31:0] inst; // @[rvdpath.scala 88:19:@3516.4]
  wire [4:0] rs1_addr; // @[rvdpath.scala 99:24:@3519.4]
  wire  _T_131; // @[rvdpath.scala 101:33:@3521.4]
  wire [31:0] _GEN_9; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_10; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_11; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_12; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_13; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_14; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_15; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_16; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_17; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_18; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_19; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_20; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_21; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_22; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_23; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_24; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_25; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_26; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_27; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_28; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_29; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_30; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_31; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_32; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_33; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_34; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_35; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_36; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_37; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_38; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] _GEN_39; // @[rvdpath.scala 101:23:@3522.4]
  wire [31:0] rs1_data; // @[rvdpath.scala 101:23:@3522.4]
  wire  _T_195; // @[Mux.scala 46:19:@3569.4]
  wire  _T_193; // @[Mux.scala 46:19:@3567.4]
  wire [31:0] z_imm; // @[Cat.scala 30:58:@3566.4]
  wire [31:0] _T_194; // @[Mux.scala 46:16:@3568.4]
  wire [31:0] _T_196; // @[Mux.scala 46:16:@3570.4]
  wire [31:0] alu_opd1; // @[Mux.scala 46:16:@3572.4]
  wire  _T_209; // @[Mux.scala 46:19:@3583.4]
  wire [4:0] rs2_addr; // @[rvdpath.scala 100:24:@3520.4]
  wire  _T_135; // @[rvdpath.scala 102:33:@3523.4]
  wire [31:0] _GEN_40; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_41; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_42; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_43; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_44; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_45; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_46; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_47; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_48; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_49; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_50; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_51; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_52; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_53; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_54; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_55; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_56; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_57; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_58; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_59; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_60; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_61; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_62; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_63; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_64; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_65; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_66; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_67; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_68; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_69; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] _GEN_70; // @[rvdpath.scala 102:23:@3524.4]
  wire [31:0] rs2_data; // @[rvdpath.scala 102:23:@3524.4]
  wire  _T_207; // @[Mux.scala 46:19:@3581.4]
  wire  _T_138; // @[rvdpath.scala 105:34:@3525.4]
  wire [19:0] _T_142; // @[Bitwise.scala 72:12:@3527.4]
  wire [11:0] _T_143; // @[rvdpath.scala 105:45:@3528.4]
  wire [31:0] i_sext; // @[Cat.scala 30:58:@3529.4]
  wire  _T_205; // @[Mux.scala 46:19:@3579.4]
  wire [6:0] _T_149; // @[rvdpath.scala 106:45:@3533.4]
  wire [26:0] _T_151; // @[Cat.scala 30:58:@3535.4]
  wire [4:0] _T_150; // @[rvdpath.scala 106:59:@3534.4]
  wire [31:0] s_sext; // @[Cat.scala 30:58:@3536.4]
  wire  _T_203; // @[Mux.scala 46:19:@3577.4]
  wire [18:0] _T_156; // @[Bitwise.scala 72:12:@3539.4]
  wire [19:0] _T_164; // @[Cat.scala 30:58:@3546.4]
  wire  _T_158; // @[rvdpath.scala 107:55:@3541.4]
  wire [20:0] _T_165; // @[Cat.scala 30:58:@3547.4]
  wire [5:0] _T_159; // @[rvdpath.scala 107:64:@3542.4]
  wire [3:0] _T_160; // @[rvdpath.scala 107:77:@3543.4]
  wire [9:0] _T_162; // @[Cat.scala 30:58:@3544.4]
  wire [10:0] _T_163; // @[Cat.scala 30:58:@3545.4]
  wire [31:0] b_sext; // @[Cat.scala 30:58:@3548.4]
  wire  _T_201; // @[Mux.scala 46:19:@3575.4]
  wire [19:0] _T_166; // @[rvdpath.scala 108:26:@3549.4]
  wire [31:0] u_sext; // @[Cat.scala 30:58:@3551.4]
  wire  _T_199; // @[Mux.scala 46:19:@3573.4]
  wire [10:0] _T_176; // @[Bitwise.scala 72:12:@3554.4]
  wire [11:0] _T_184; // @[Cat.scala 30:58:@3561.4]
  wire [7:0] _T_178; // @[rvdpath.scala 109:55:@3556.4]
  wire [19:0] _T_185; // @[Cat.scala 30:58:@3562.4]
  wire  _T_179; // @[rvdpath.scala 109:68:@3557.4]
  wire [9:0] _T_180; // @[rvdpath.scala 109:78:@3558.4]
  wire [10:0] _T_182; // @[Cat.scala 30:58:@3559.4]
  wire [11:0] _T_183; // @[Cat.scala 30:58:@3560.4]
  wire [31:0] j_sext; // @[Cat.scala 30:58:@3563.4]
  wire [31:0] _T_200; // @[Mux.scala 46:16:@3574.4]
  wire [31:0] _T_202; // @[Mux.scala 46:16:@3576.4]
  wire [31:0] _T_204; // @[Mux.scala 46:16:@3578.4]
  wire [31:0] _T_206; // @[Mux.scala 46:16:@3580.4]
  wire [31:0] _T_208; // @[Mux.scala 46:16:@3582.4]
  wire [31:0] alu_opd2; // @[Mux.scala 46:16:@3584.4]
  wire [32:0] _T_219; // @[rvdpath.scala 153:38:@3596.4]
  wire [31:0] _T_220; // @[rvdpath.scala 153:38:@3597.4]
  wire  _T_259; // @[Mux.scala 46:19:@3636.4]
  wire [32:0] _T_221; // @[rvdpath.scala 154:38:@3598.4]
  wire [32:0] _T_222; // @[rvdpath.scala 154:38:@3599.4]
  wire [31:0] _T_223; // @[rvdpath.scala 154:38:@3600.4]
  wire  _T_257; // @[Mux.scala 46:19:@3634.4]
  wire [4:0] _T_224; // @[rvdpath.scala 158:49:@3601.4]
  wire [62:0] _GEN_489; // @[rvdpath.scala 158:38:@3602.4]
  wire [62:0] _T_225; // @[rvdpath.scala 158:38:@3602.4]
  wire  _T_255; // @[Mux.scala 46:19:@3632.4]
  wire [31:0] _T_226; // @[rvdpath.scala 159:38:@3603.4]
  wire [31:0] _T_227; // @[rvdpath.scala 159:56:@3604.4]
  wire  _T_228; // @[rvdpath.scala 159:45:@3605.4]
  wire  _T_253; // @[Mux.scala 46:19:@3630.4]
  wire  _T_229; // @[rvdpath.scala 160:38:@3606.4]
  wire  _T_251; // @[Mux.scala 46:19:@3628.4]
  wire [31:0] _T_230; // @[rvdpath.scala 161:38:@3607.4]
  wire  _T_249; // @[Mux.scala 46:19:@3626.4]
  wire [31:0] _T_232; // @[rvdpath.scala 162:38:@3609.4]
  wire  _T_247; // @[Mux.scala 46:19:@3624.4]
  wire [31:0] _T_235; // @[rvdpath.scala 163:45:@3612.4]
  wire [31:0] _T_236; // @[rvdpath.scala 163:78:@3613.4]
  wire  _T_245; // @[Mux.scala 46:19:@3622.4]
  wire [31:0] _T_237; // @[rvdpath.scala 164:38:@3614.4]
  wire  _T_243; // @[Mux.scala 46:19:@3620.4]
  wire [31:0] _T_238; // @[rvdpath.scala 165:38:@3615.4]
  wire  _T_241; // @[Mux.scala 46:19:@3618.4]
  wire  _T_239; // @[Mux.scala 46:19:@3616.4]
  wire [31:0] _T_240; // @[Mux.scala 46:16:@3617.4]
  wire [31:0] _T_242; // @[Mux.scala 46:16:@3619.4]
  wire [31:0] _T_244; // @[Mux.scala 46:16:@3621.4]
  wire [31:0] _T_246; // @[Mux.scala 46:16:@3623.4]
  wire [31:0] _T_248; // @[Mux.scala 46:16:@3625.4]
  wire [31:0] _T_250; // @[Mux.scala 46:16:@3627.4]
  wire [31:0] _T_252; // @[Mux.scala 46:16:@3629.4]
  wire [31:0] _T_254; // @[Mux.scala 46:16:@3631.4]
  wire [31:0] _T_256; // @[Mux.scala 46:16:@3633.4]
  wire [62:0] _T_258; // @[Mux.scala 46:16:@3635.4]
  wire [62:0] _T_260; // @[Mux.scala 46:16:@3637.4]
  wire [62:0] _T_262; // @[Mux.scala 46:16:@3639.4]
  wire [31:0] alu_out; // @[rvdpath.scala 169:6:@3640.4]
  wire [31:0] _T_76; // @[Mux.scala 46:16:@3492.4]
  wire  _T_77; // @[Mux.scala 46:19:@3493.4]
  wire  _T_285; // @[Mux.scala 46:19:@3660.4]
  wire  bcmp_eq; // @[rvdpath.scala 140:26:@3588.4]
  wire [31:0] _T_263; // @[rvdpath.scala 177:35:@3641.4]
  wire  _T_283; // @[Mux.scala 46:19:@3658.4]
  wire  _T_265; // @[rvdpath.scala 178:36:@3642.4]
  wire [31:0] _T_266; // @[rvdpath.scala 178:35:@3643.4]
  wire  _T_281; // @[Mux.scala 46:19:@3656.4]
  wire [31:0] _T_214; // @[rvdpath.scala 141:26:@3590.4]
  wire [31:0] _T_215; // @[rvdpath.scala 141:44:@3591.4]
  wire  bcmp_lt; // @[rvdpath.scala 141:33:@3592.4]
  wire [31:0] _T_267; // @[rvdpath.scala 179:35:@3644.4]
  wire  _T_279; // @[Mux.scala 46:19:@3654.4]
  wire  _T_269; // @[rvdpath.scala 180:36:@3645.4]
  wire [31:0] _T_270; // @[rvdpath.scala 180:35:@3646.4]
  wire  _T_277; // @[Mux.scala 46:19:@3652.4]
  wire  bcmp_ltu; // @[rvdpath.scala 142:34:@3594.4]
  wire [31:0] _T_271; // @[rvdpath.scala 181:36:@3647.4]
  wire  _T_275; // @[Mux.scala 46:19:@3650.4]
  wire  _T_273; // @[rvdpath.scala 182:37:@3648.4]
  wire [31:0] _T_274; // @[rvdpath.scala 182:36:@3649.4]
  wire [31:0] _T_276; // @[Mux.scala 46:16:@3651.4]
  wire [31:0] _T_278; // @[Mux.scala 46:16:@3653.4]
  wire [31:0] _T_280; // @[Mux.scala 46:16:@3655.4]
  wire [31:0] _T_282; // @[Mux.scala 46:16:@3657.4]
  wire [31:0] _T_284; // @[Mux.scala 46:16:@3659.4]
  wire [31:0] pc_br; // @[Mux.scala 46:16:@3661.4]
  wire [31:0] _T_78; // @[Mux.scala 46:16:@3494.4]
  wire  _T_79; // @[Mux.scala 46:19:@3495.4]
  wire [31:0] pc_next; // @[Mux.scala 46:16:@3496.4]
  wire  _T_84; // @[rvdpath.scala 77:42:@3504.4]
  wire  _T_85; // @[rvdpath.scala 77:40:@3505.4]
  wire  _T_86; // @[rvdpath.scala 78:39:@3506.4]
  wire  _T_87; // @[rvdpath.scala 78:51:@3507.4]
  wire  _T_88; // @[rvdpath.scala 77:63:@3508.4]
  wire  _T_90; // @[rvdpath.scala 79:41:@3509.4]
  wire  _T_91; // @[rvdpath.scala 79:39:@3510.4]
  wire  _T_92; // @[rvdpath.scala 79:52:@3511.4]
  wire  pc_update; // @[rvdpath.scala 78:73:@3512.4]
  wire [31:0] _GEN_8; // @[rvdpath.scala 81:21:@3513.4]
  wire  _T_291; // @[Mux.scala 46:19:@3671.4]
  wire [1:0] _T_292; // @[Mux.scala 46:16:@3672.4]
  wire  _T_293; // @[Mux.scala 46:19:@3673.4]
  wire [1:0] _T_294; // @[Mux.scala 46:16:@3674.4]
  wire  _T_295; // @[Mux.scala 46:19:@3675.4]
  wire [1:0] _T_296; // @[Mux.scala 46:16:@3676.4]
  wire  _T_297; // @[Mux.scala 46:19:@3677.4]
  wire [1:0] _T_298; // @[Mux.scala 46:16:@3678.4]
  wire  _T_299; // @[Mux.scala 46:19:@3679.4]
  wire [1:0] mem_type; // @[Mux.scala 46:16:@3680.4]
  wire  _T_301; // @[Conditional.scala 37:30:@3685.6]
  wire  _T_304; // @[rvdpath.scala 220:49:@3687.8]
  wire [31:0] _T_306; // @[rvdpath.scala 220:40:@3688.8]
  wire [31:0] _GEN_71; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_72; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_73; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_74; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_75; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_76; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_77; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_78; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_79; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_80; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_81; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_82; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_83; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_84; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_85; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_86; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_87; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_88; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_89; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_90; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_91; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_92; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_93; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_94; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_95; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_96; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_97; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_98; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_99; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_100; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_101; // @[rvdpath.scala 220:34:@3689.8]
  wire [31:0] _GEN_102; // @[rvdpath.scala 220:34:@3689.8]
  wire  _T_307; // @[Conditional.scala 37:30:@3692.8]
  wire  _T_309; // @[rvdpath.scala 228:77:@3695.12]
  wire [23:0] _T_313; // @[Bitwise.scala 72:12:@3697.12]
  wire [7:0] _T_314; // @[rvdpath.scala 228:100:@3698.12]
  wire [31:0] _T_315; // @[Cat.scala 30:58:@3699.12]
  wire  _T_316; // @[rvdpath.scala 229:77:@3700.12]
  wire [15:0] _T_320; // @[Bitwise.scala 72:12:@3702.12]
  wire [15:0] _T_321; // @[rvdpath.scala 229:101:@3703.12]
  wire [31:0] _T_322; // @[Cat.scala 30:58:@3704.12]
  wire [31:0] _T_329; // @[Cat.scala 30:58:@3707.12]
  wire [31:0] _T_336; // @[Cat.scala 30:58:@3710.12]
  wire [31:0] _T_338; // @[Mux.scala 46:16:@3712.12]
  wire [31:0] _T_340; // @[Mux.scala 46:16:@3714.12]
  wire [31:0] _T_342; // @[Mux.scala 46:16:@3716.12]
  wire [31:0] _T_344; // @[Mux.scala 46:16:@3718.12]
  wire [31:0] _T_346; // @[Mux.scala 46:16:@3720.12]
  wire [31:0] _T_351; // @[rvdpath.scala 236:44:@3722.12]
  wire [31:0] _GEN_103; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_104; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_105; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_106; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_107; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_108; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_109; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_110; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_111; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_112; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_113; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_114; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_115; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_116; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_117; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_118; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_119; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_120; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_121; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_122; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_123; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_124; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_125; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_126; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_127; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_128; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_129; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_130; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_131; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_132; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_133; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_134; // @[rvdpath.scala 236:38:@3723.12]
  wire [31:0] _GEN_135; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_136; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_137; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_138; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_139; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_140; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_141; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_142; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_143; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_144; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_145; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_146; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_147; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_148; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_149; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_150; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_151; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_152; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_153; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_154; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_155; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_156; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_157; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_158; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_159; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_160; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_161; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_162; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_163; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_164; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_165; // @[rvdpath.scala 223:42:@3694.10]
  wire [31:0] _GEN_166; // @[rvdpath.scala 223:42:@3694.10]
  wire  _T_352; // @[Conditional.scala 37:30:@3727.10]
  wire [31:0] _T_357; // @[rvdpath.scala 241:40:@3730.12]
  wire [31:0] _GEN_167; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_168; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_169; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_170; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_171; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_172; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_173; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_174; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_175; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_176; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_177; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_178; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_179; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_180; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_181; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_182; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_183; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_184; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_185; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_186; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_187; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_188; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_189; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_190; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_191; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_192; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_193; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_194; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_195; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_196; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_197; // @[rvdpath.scala 241:34:@3731.12]
  wire [31:0] _GEN_198; // @[rvdpath.scala 241:34:@3731.12]
  wire  _T_358; // @[Conditional.scala 37:30:@3734.12]
  wire [31:0] csr_rdata; // @[rvdpath.scala 192:25:@3664.4]
  wire [31:0] _T_363; // @[rvdpath.scala 245:40:@3737.14]
  wire [31:0] _GEN_199; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_200; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_201; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_202; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_203; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_204; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_205; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_206; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_207; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_208; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_209; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_210; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_211; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_212; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_213; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_214; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_215; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_216; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_217; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_218; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_219; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_220; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_221; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_222; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_223; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_224; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_225; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_226; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_227; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_228; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_229; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_230; // @[rvdpath.scala 245:34:@3738.14]
  wire [31:0] _GEN_231; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_232; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_233; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_234; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_235; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_236; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_237; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_238; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_239; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_240; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_241; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_242; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_243; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_244; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_245; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_246; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_247; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_248; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_249; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_250; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_251; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_252; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_253; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_254; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_255; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_256; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_257; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_258; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_259; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_260; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_261; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_262; // @[Conditional.scala 39:67:@3735.12]
  wire [31:0] _GEN_263; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_264; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_265; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_266; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_267; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_268; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_269; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_270; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_271; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_272; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_273; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_274; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_275; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_276; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_277; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_278; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_279; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_280; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_281; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_282; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_283; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_284; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_285; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_286; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_287; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_288; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_289; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_290; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_291; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_292; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_293; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_294; // @[Conditional.scala 39:67:@3728.10]
  wire [31:0] _GEN_295; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_296; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_297; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_298; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_299; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_300; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_301; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_302; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_303; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_304; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_305; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_306; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_307; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_308; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_309; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_310; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_311; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_312; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_313; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_314; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_315; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_316; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_317; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_318; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_319; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_320; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_321; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_322; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_323; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_324; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_325; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_326; // @[Conditional.scala 39:67:@3693.8]
  wire [31:0] _GEN_327; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_328; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_329; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_330; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_331; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_332; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_333; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_334; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_335; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_336; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_337; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_338; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_339; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_340; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_341; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_342; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_343; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_344; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_345; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_346; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_347; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_348; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_349; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_350; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_351; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_352; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_353; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_354; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_355; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_356; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_357; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_358; // @[Conditional.scala 40:58:@3686.6]
  wire [31:0] _GEN_359; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_360; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_361; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_362; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_363; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_364; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_365; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_366; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_367; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_368; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_369; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_370; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_371; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_372; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_373; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_374; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_375; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_376; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_377; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_378; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_379; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_380; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_381; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_382; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_383; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_384; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_385; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_386; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_387; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_388; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_389; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_390; // @[rvdpath.scala 216:47:@3684.4]
  wire [31:0] _GEN_391; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_392; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_393; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_394; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_395; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_396; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_397; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_398; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_399; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_400; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_401; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_402; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_403; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_404; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_405; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_406; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_407; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_408; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_409; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_410; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_411; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_412; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_413; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_414; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_415; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_416; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_417; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_418; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_419; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_420; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_421; // @[rvdpath.scala 265:21:@3755.4]
  wire [31:0] _GEN_422; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_423; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_424; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_425; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_426; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_427; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_428; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_429; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_430; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_431; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_432; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_433; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_434; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_435; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_436; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_437; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_438; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_439; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_440; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_441; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_442; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_443; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_444; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_445; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_446; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_447; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_448; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_449; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_450; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_451; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_452; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_453; // @[rvdpath.scala 267:33:@3757.6]
  wire [31:0] _GEN_454; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_455; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_456; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_457; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_458; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_459; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_460; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_461; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_462; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_463; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_464; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_465; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_466; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_467; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_468; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_469; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_470; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_471; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_472; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_473; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_474; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_475; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_476; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_477; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_478; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_479; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_480; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_481; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_482; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_483; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_484; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_485; // @[rvdpath.scala 266:26:@3756.4]
  wire [31:0] _GEN_486; // @[rvdpath.scala 271:26:@3760.4]
  wire  _GEN_487; // @[rvdpath.scala 271:26:@3760.4]
  wire  _GEN_488; // @[rvdpath.scala 271:26:@3760.4]
  rvcsr csr ( // @[rvdpath.scala 251:21:@3741.4]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_addr(csr_io_addr),
    .io_wdata(csr_io_wdata),
    .io_rdata(csr_io_rdata),
    .io_op(csr_io_op),
    .io_core_pc(csr_io_core_pc),
    .io_core_excp(csr_io_core_excp),
    .io_core_cause(csr_io_core_cause),
    .io_csr_excp(csr_io_csr_excp),
    .io_csr_evec(csr_io_csr_evec)
  );
  assign _T_71 = pc + 32'h4; // @[rvdpath.scala 52:17:@3486.4]
  assign pc_a4 = _T_71[31:0]; // @[rvdpath.scala 52:17:@3487.4]
  assign _T_73 = 2'h3 == io_c2d_pc_sel; // @[Mux.scala 46:19:@3489.4]
  assign pc_ex = csr_io_csr_evec; // @[rvdpath.scala 50:21:@3485.4]
  assign _T_74 = _T_73 ? pc_ex : pc_a4; // @[Mux.scala 46:16:@3490.4]
  assign _T_75 = 2'h2 == io_c2d_pc_sel; // @[Mux.scala 46:19:@3491.4]
  assign _T_261 = 4'h0 == io_c2d_alu_func; // @[Mux.scala 46:19:@3638.4]
  assign _T_197 = 2'h0 == io_c2d_op1_sel; // @[Mux.scala 46:19:@3571.4]
  assign inst = io_imem_resp_valid ? io_imem_resp_data : 32'h13; // @[rvdpath.scala 88:19:@3516.4]
  assign rs1_addr = inst[19:15]; // @[rvdpath.scala 99:24:@3519.4]
  assign _T_131 = rs1_addr != 5'h0; // @[rvdpath.scala 101:33:@3521.4]
  assign _GEN_9 = 5'h1 == rs1_addr ? regfile_1 : regfile_0; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_10 = 5'h2 == rs1_addr ? regfile_2 : _GEN_9; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_11 = 5'h3 == rs1_addr ? regfile_3 : _GEN_10; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_12 = 5'h4 == rs1_addr ? regfile_4 : _GEN_11; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_13 = 5'h5 == rs1_addr ? regfile_5 : _GEN_12; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_14 = 5'h6 == rs1_addr ? regfile_6 : _GEN_13; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_15 = 5'h7 == rs1_addr ? regfile_7 : _GEN_14; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_16 = 5'h8 == rs1_addr ? regfile_8 : _GEN_15; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_17 = 5'h9 == rs1_addr ? regfile_9 : _GEN_16; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_18 = 5'ha == rs1_addr ? regfile_10 : _GEN_17; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_19 = 5'hb == rs1_addr ? regfile_11 : _GEN_18; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_20 = 5'hc == rs1_addr ? regfile_12 : _GEN_19; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_21 = 5'hd == rs1_addr ? regfile_13 : _GEN_20; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_22 = 5'he == rs1_addr ? regfile_14 : _GEN_21; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_23 = 5'hf == rs1_addr ? regfile_15 : _GEN_22; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_24 = 5'h10 == rs1_addr ? regfile_16 : _GEN_23; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_25 = 5'h11 == rs1_addr ? regfile_17 : _GEN_24; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_26 = 5'h12 == rs1_addr ? regfile_18 : _GEN_25; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_27 = 5'h13 == rs1_addr ? regfile_19 : _GEN_26; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_28 = 5'h14 == rs1_addr ? regfile_20 : _GEN_27; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_29 = 5'h15 == rs1_addr ? regfile_21 : _GEN_28; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_30 = 5'h16 == rs1_addr ? regfile_22 : _GEN_29; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_31 = 5'h17 == rs1_addr ? regfile_23 : _GEN_30; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_32 = 5'h18 == rs1_addr ? regfile_24 : _GEN_31; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_33 = 5'h19 == rs1_addr ? regfile_25 : _GEN_32; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_34 = 5'h1a == rs1_addr ? regfile_26 : _GEN_33; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_35 = 5'h1b == rs1_addr ? regfile_27 : _GEN_34; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_36 = 5'h1c == rs1_addr ? regfile_28 : _GEN_35; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_37 = 5'h1d == rs1_addr ? regfile_29 : _GEN_36; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_38 = 5'h1e == rs1_addr ? regfile_30 : _GEN_37; // @[rvdpath.scala 101:23:@3522.4]
  assign _GEN_39 = 5'h1f == rs1_addr ? regfile_31 : _GEN_38; // @[rvdpath.scala 101:23:@3522.4]
  assign rs1_data = _T_131 ? _GEN_39 : 32'h0; // @[rvdpath.scala 101:23:@3522.4]
  assign _T_195 = 2'h1 == io_c2d_op1_sel; // @[Mux.scala 46:19:@3569.4]
  assign _T_193 = 2'h2 == io_c2d_op1_sel; // @[Mux.scala 46:19:@3567.4]
  assign z_imm = {27'h0,rs1_addr}; // @[Cat.scala 30:58:@3566.4]
  assign _T_194 = _T_193 ? z_imm : 32'h0; // @[Mux.scala 46:16:@3568.4]
  assign _T_196 = _T_195 ? pc : _T_194; // @[Mux.scala 46:16:@3570.4]
  assign alu_opd1 = _T_197 ? rs1_data : _T_196; // @[Mux.scala 46:16:@3572.4]
  assign _T_209 = 3'h0 == io_c2d_op2_sel; // @[Mux.scala 46:19:@3583.4]
  assign rs2_addr = inst[24:20]; // @[rvdpath.scala 100:24:@3520.4]
  assign _T_135 = rs2_addr != 5'h0; // @[rvdpath.scala 102:33:@3523.4]
  assign _GEN_40 = 5'h1 == rs2_addr ? regfile_1 : regfile_0; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_41 = 5'h2 == rs2_addr ? regfile_2 : _GEN_40; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_42 = 5'h3 == rs2_addr ? regfile_3 : _GEN_41; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_43 = 5'h4 == rs2_addr ? regfile_4 : _GEN_42; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_44 = 5'h5 == rs2_addr ? regfile_5 : _GEN_43; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_45 = 5'h6 == rs2_addr ? regfile_6 : _GEN_44; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_46 = 5'h7 == rs2_addr ? regfile_7 : _GEN_45; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_47 = 5'h8 == rs2_addr ? regfile_8 : _GEN_46; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_48 = 5'h9 == rs2_addr ? regfile_9 : _GEN_47; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_49 = 5'ha == rs2_addr ? regfile_10 : _GEN_48; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_50 = 5'hb == rs2_addr ? regfile_11 : _GEN_49; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_51 = 5'hc == rs2_addr ? regfile_12 : _GEN_50; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_52 = 5'hd == rs2_addr ? regfile_13 : _GEN_51; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_53 = 5'he == rs2_addr ? regfile_14 : _GEN_52; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_54 = 5'hf == rs2_addr ? regfile_15 : _GEN_53; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_55 = 5'h10 == rs2_addr ? regfile_16 : _GEN_54; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_56 = 5'h11 == rs2_addr ? regfile_17 : _GEN_55; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_57 = 5'h12 == rs2_addr ? regfile_18 : _GEN_56; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_58 = 5'h13 == rs2_addr ? regfile_19 : _GEN_57; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_59 = 5'h14 == rs2_addr ? regfile_20 : _GEN_58; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_60 = 5'h15 == rs2_addr ? regfile_21 : _GEN_59; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_61 = 5'h16 == rs2_addr ? regfile_22 : _GEN_60; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_62 = 5'h17 == rs2_addr ? regfile_23 : _GEN_61; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_63 = 5'h18 == rs2_addr ? regfile_24 : _GEN_62; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_64 = 5'h19 == rs2_addr ? regfile_25 : _GEN_63; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_65 = 5'h1a == rs2_addr ? regfile_26 : _GEN_64; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_66 = 5'h1b == rs2_addr ? regfile_27 : _GEN_65; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_67 = 5'h1c == rs2_addr ? regfile_28 : _GEN_66; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_68 = 5'h1d == rs2_addr ? regfile_29 : _GEN_67; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_69 = 5'h1e == rs2_addr ? regfile_30 : _GEN_68; // @[rvdpath.scala 102:23:@3524.4]
  assign _GEN_70 = 5'h1f == rs2_addr ? regfile_31 : _GEN_69; // @[rvdpath.scala 102:23:@3524.4]
  assign rs2_data = _T_135 ? _GEN_70 : 32'h0; // @[rvdpath.scala 102:23:@3524.4]
  assign _T_207 = 3'h1 == io_c2d_op2_sel; // @[Mux.scala 46:19:@3581.4]
  assign _T_138 = inst[31]; // @[rvdpath.scala 105:34:@3525.4]
  assign _T_142 = _T_138 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@3527.4]
  assign _T_143 = inst[31:20]; // @[rvdpath.scala 105:45:@3528.4]
  assign i_sext = {_T_142,_T_143}; // @[Cat.scala 30:58:@3529.4]
  assign _T_205 = 3'h2 == io_c2d_op2_sel; // @[Mux.scala 46:19:@3579.4]
  assign _T_149 = inst[31:25]; // @[rvdpath.scala 106:45:@3533.4]
  assign _T_151 = {_T_142,_T_149}; // @[Cat.scala 30:58:@3535.4]
  assign _T_150 = inst[11:7]; // @[rvdpath.scala 106:59:@3534.4]
  assign s_sext = {_T_151,_T_150}; // @[Cat.scala 30:58:@3536.4]
  assign _T_203 = 3'h3 == io_c2d_op2_sel; // @[Mux.scala 46:19:@3577.4]
  assign _T_156 = _T_138 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12:@3539.4]
  assign _T_164 = {_T_156,_T_138}; // @[Cat.scala 30:58:@3546.4]
  assign _T_158 = inst[7]; // @[rvdpath.scala 107:55:@3541.4]
  assign _T_165 = {_T_164,_T_158}; // @[Cat.scala 30:58:@3547.4]
  assign _T_159 = inst[30:25]; // @[rvdpath.scala 107:64:@3542.4]
  assign _T_160 = inst[11:8]; // @[rvdpath.scala 107:77:@3543.4]
  assign _T_162 = {_T_159,_T_160}; // @[Cat.scala 30:58:@3544.4]
  assign _T_163 = {_T_162,1'h0}; // @[Cat.scala 30:58:@3545.4]
  assign b_sext = {_T_165,_T_163}; // @[Cat.scala 30:58:@3548.4]
  assign _T_201 = 3'h4 == io_c2d_op2_sel; // @[Mux.scala 46:19:@3575.4]
  assign _T_166 = inst[31:12]; // @[rvdpath.scala 108:26:@3549.4]
  assign u_sext = {_T_166,12'h0}; // @[Cat.scala 30:58:@3551.4]
  assign _T_199 = 3'h5 == io_c2d_op2_sel; // @[Mux.scala 46:19:@3573.4]
  assign _T_176 = _T_138 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12:@3554.4]
  assign _T_184 = {_T_176,_T_138}; // @[Cat.scala 30:58:@3561.4]
  assign _T_178 = inst[19:12]; // @[rvdpath.scala 109:55:@3556.4]
  assign _T_185 = {_T_184,_T_178}; // @[Cat.scala 30:58:@3562.4]
  assign _T_179 = inst[20]; // @[rvdpath.scala 109:68:@3557.4]
  assign _T_180 = inst[30:21]; // @[rvdpath.scala 109:78:@3558.4]
  assign _T_182 = {_T_179,_T_180}; // @[Cat.scala 30:58:@3559.4]
  assign _T_183 = {_T_182,1'h0}; // @[Cat.scala 30:58:@3560.4]
  assign j_sext = {_T_185,_T_183}; // @[Cat.scala 30:58:@3563.4]
  assign _T_200 = _T_199 ? j_sext : 32'h0; // @[Mux.scala 46:16:@3574.4]
  assign _T_202 = _T_201 ? u_sext : _T_200; // @[Mux.scala 46:16:@3576.4]
  assign _T_204 = _T_203 ? b_sext : _T_202; // @[Mux.scala 46:16:@3578.4]
  assign _T_206 = _T_205 ? s_sext : _T_204; // @[Mux.scala 46:16:@3580.4]
  assign _T_208 = _T_207 ? i_sext : _T_206; // @[Mux.scala 46:16:@3582.4]
  assign alu_opd2 = _T_209 ? rs2_data : _T_208; // @[Mux.scala 46:16:@3584.4]
  assign _T_219 = alu_opd1 + alu_opd2; // @[rvdpath.scala 153:38:@3596.4]
  assign _T_220 = _T_219[31:0]; // @[rvdpath.scala 153:38:@3597.4]
  assign _T_259 = 4'h8 == io_c2d_alu_func; // @[Mux.scala 46:19:@3636.4]
  assign _T_221 = alu_opd1 - alu_opd2; // @[rvdpath.scala 154:38:@3598.4]
  assign _T_222 = $unsigned(_T_221); // @[rvdpath.scala 154:38:@3599.4]
  assign _T_223 = _T_222[31:0]; // @[rvdpath.scala 154:38:@3600.4]
  assign _T_257 = 4'h1 == io_c2d_alu_func; // @[Mux.scala 46:19:@3634.4]
  assign _T_224 = alu_opd2[4:0]; // @[rvdpath.scala 158:49:@3601.4]
  assign _GEN_489 = {{31'd0}, alu_opd1}; // @[rvdpath.scala 158:38:@3602.4]
  assign _T_225 = _GEN_489 << _T_224; // @[rvdpath.scala 158:38:@3602.4]
  assign _T_255 = 4'h2 == io_c2d_alu_func; // @[Mux.scala 46:19:@3632.4]
  assign _T_226 = $signed(alu_opd1); // @[rvdpath.scala 159:38:@3603.4]
  assign _T_227 = $signed(alu_opd2); // @[rvdpath.scala 159:56:@3604.4]
  assign _T_228 = $signed(_T_226) < $signed(_T_227); // @[rvdpath.scala 159:45:@3605.4]
  assign _T_253 = 4'h3 == io_c2d_alu_func; // @[Mux.scala 46:19:@3630.4]
  assign _T_229 = alu_opd1 < alu_opd2; // @[rvdpath.scala 160:38:@3606.4]
  assign _T_251 = 4'h4 == io_c2d_alu_func; // @[Mux.scala 46:19:@3628.4]
  assign _T_230 = alu_opd1 ^ alu_opd2; // @[rvdpath.scala 161:38:@3607.4]
  assign _T_249 = 4'h5 == io_c2d_alu_func; // @[Mux.scala 46:19:@3626.4]
  assign _T_232 = alu_opd1 >> _T_224; // @[rvdpath.scala 162:38:@3609.4]
  assign _T_247 = 4'hd == io_c2d_alu_func; // @[Mux.scala 46:19:@3624.4]
  assign _T_235 = $signed(_T_226) >>> _T_224; // @[rvdpath.scala 163:45:@3612.4]
  assign _T_236 = $unsigned(_T_235); // @[rvdpath.scala 163:78:@3613.4]
  assign _T_245 = 4'h6 == io_c2d_alu_func; // @[Mux.scala 46:19:@3622.4]
  assign _T_237 = alu_opd1 | alu_opd2; // @[rvdpath.scala 164:38:@3614.4]
  assign _T_243 = 4'h7 == io_c2d_alu_func; // @[Mux.scala 46:19:@3620.4]
  assign _T_238 = alu_opd1 & alu_opd2; // @[rvdpath.scala 165:38:@3615.4]
  assign _T_241 = 4'ha == io_c2d_alu_func; // @[Mux.scala 46:19:@3618.4]
  assign _T_239 = 4'hb == io_c2d_alu_func; // @[Mux.scala 46:19:@3616.4]
  assign _T_240 = _T_239 ? alu_opd2 : 32'h0; // @[Mux.scala 46:16:@3617.4]
  assign _T_242 = _T_241 ? alu_opd1 : _T_240; // @[Mux.scala 46:16:@3619.4]
  assign _T_244 = _T_243 ? _T_238 : _T_242; // @[Mux.scala 46:16:@3621.4]
  assign _T_246 = _T_245 ? _T_237 : _T_244; // @[Mux.scala 46:16:@3623.4]
  assign _T_248 = _T_247 ? _T_236 : _T_246; // @[Mux.scala 46:16:@3625.4]
  assign _T_250 = _T_249 ? _T_232 : _T_248; // @[Mux.scala 46:16:@3627.4]
  assign _T_252 = _T_251 ? _T_230 : _T_250; // @[Mux.scala 46:16:@3629.4]
  assign _T_254 = _T_253 ? {{31'd0}, _T_229} : _T_252; // @[Mux.scala 46:16:@3631.4]
  assign _T_256 = _T_255 ? {{31'd0}, _T_228} : _T_254; // @[Mux.scala 46:16:@3633.4]
  assign _T_258 = _T_257 ? _T_225 : {{31'd0}, _T_256}; // @[Mux.scala 46:16:@3635.4]
  assign _T_260 = _T_259 ? {{31'd0}, _T_223} : _T_258; // @[Mux.scala 46:16:@3637.4]
  assign _T_262 = _T_261 ? {{31'd0}, _T_220} : _T_260; // @[Mux.scala 46:16:@3639.4]
  assign alu_out = _T_262[31:0]; // @[rvdpath.scala 169:6:@3640.4]
  assign _T_76 = _T_75 ? alu_out : _T_74; // @[Mux.scala 46:16:@3492.4]
  assign _T_77 = 2'h1 == io_c2d_pc_sel; // @[Mux.scala 46:19:@3493.4]
  assign _T_285 = 3'h0 == io_c2d_br_sel; // @[Mux.scala 46:19:@3660.4]
  assign bcmp_eq = rs1_data == rs2_data; // @[rvdpath.scala 140:26:@3588.4]
  assign _T_263 = bcmp_eq ? alu_out : pc_a4; // @[rvdpath.scala 177:35:@3641.4]
  assign _T_283 = 3'h1 == io_c2d_br_sel; // @[Mux.scala 46:19:@3658.4]
  assign _T_265 = bcmp_eq == 1'h0; // @[rvdpath.scala 178:36:@3642.4]
  assign _T_266 = _T_265 ? alu_out : pc_a4; // @[rvdpath.scala 178:35:@3643.4]
  assign _T_281 = 3'h2 == io_c2d_br_sel; // @[Mux.scala 46:19:@3656.4]
  assign _T_214 = $signed(rs1_data); // @[rvdpath.scala 141:26:@3590.4]
  assign _T_215 = $signed(rs2_data); // @[rvdpath.scala 141:44:@3591.4]
  assign bcmp_lt = $signed(_T_214) < $signed(_T_215); // @[rvdpath.scala 141:33:@3592.4]
  assign _T_267 = bcmp_lt ? alu_out : pc_a4; // @[rvdpath.scala 179:35:@3644.4]
  assign _T_279 = 3'h3 == io_c2d_br_sel; // @[Mux.scala 46:19:@3654.4]
  assign _T_269 = bcmp_lt == 1'h0; // @[rvdpath.scala 180:36:@3645.4]
  assign _T_270 = _T_269 ? alu_out : pc_a4; // @[rvdpath.scala 180:35:@3646.4]
  assign _T_277 = 3'h4 == io_c2d_br_sel; // @[Mux.scala 46:19:@3652.4]
  assign bcmp_ltu = rs1_data < rs2_data; // @[rvdpath.scala 142:34:@3594.4]
  assign _T_271 = bcmp_ltu ? alu_out : pc_a4; // @[rvdpath.scala 181:36:@3647.4]
  assign _T_275 = 3'h5 == io_c2d_br_sel; // @[Mux.scala 46:19:@3650.4]
  assign _T_273 = bcmp_ltu == 1'h0; // @[rvdpath.scala 182:37:@3648.4]
  assign _T_274 = _T_273 ? alu_out : pc_a4; // @[rvdpath.scala 182:36:@3649.4]
  assign _T_276 = _T_275 ? _T_274 : pc_a4; // @[Mux.scala 46:16:@3651.4]
  assign _T_278 = _T_277 ? _T_271 : _T_276; // @[Mux.scala 46:16:@3653.4]
  assign _T_280 = _T_279 ? _T_270 : _T_278; // @[Mux.scala 46:16:@3655.4]
  assign _T_282 = _T_281 ? _T_267 : _T_280; // @[Mux.scala 46:16:@3657.4]
  assign _T_284 = _T_283 ? _T_266 : _T_282; // @[Mux.scala 46:16:@3659.4]
  assign pc_br = _T_285 ? _T_263 : _T_284; // @[Mux.scala 46:16:@3661.4]
  assign _T_78 = _T_77 ? pc_br : _T_76; // @[Mux.scala 46:16:@3494.4]
  assign _T_79 = 2'h0 == io_c2d_pc_sel; // @[Mux.scala 46:19:@3495.4]
  assign pc_next = _T_79 ? pc_a4 : _T_78; // @[Mux.scala 46:16:@3496.4]
  assign _T_84 = io_dmem_req_valid == 1'h0; // @[rvdpath.scala 77:42:@3504.4]
  assign _T_85 = io_imem_resp_valid & _T_84; // @[rvdpath.scala 77:40:@3505.4]
  assign _T_86 = io_dmem_req_valid & io_c2d_mem_wren; // @[rvdpath.scala 78:39:@3506.4]
  assign _T_87 = _T_86 & io_dmem_req_ready; // @[rvdpath.scala 78:51:@3507.4]
  assign _T_88 = _T_85 | _T_87; // @[rvdpath.scala 77:63:@3508.4]
  assign _T_90 = io_c2d_mem_wren == 1'h0; // @[rvdpath.scala 79:41:@3509.4]
  assign _T_91 = io_dmem_req_valid & _T_90; // @[rvdpath.scala 79:39:@3510.4]
  assign _T_92 = _T_91 & io_dmem_resp_valid; // @[rvdpath.scala 79:52:@3511.4]
  assign pc_update = _T_88 | _T_92; // @[rvdpath.scala 78:73:@3512.4]
  assign _GEN_8 = pc_update ? pc_next : pc; // @[rvdpath.scala 81:21:@3513.4]
  assign _T_291 = 3'h5 == io_c2d_mem_type; // @[Mux.scala 46:19:@3671.4]
  assign _T_292 = _T_291 ? 2'h2 : 2'h0; // @[Mux.scala 46:16:@3672.4]
  assign _T_293 = 3'h4 == io_c2d_mem_type; // @[Mux.scala 46:19:@3673.4]
  assign _T_294 = _T_293 ? 2'h1 : _T_292; // @[Mux.scala 46:16:@3674.4]
  assign _T_295 = 3'h2 == io_c2d_mem_type; // @[Mux.scala 46:19:@3675.4]
  assign _T_296 = _T_295 ? 2'h3 : _T_294; // @[Mux.scala 46:16:@3676.4]
  assign _T_297 = 3'h1 == io_c2d_mem_type; // @[Mux.scala 46:19:@3677.4]
  assign _T_298 = _T_297 ? 2'h2 : _T_296; // @[Mux.scala 46:16:@3678.4]
  assign _T_299 = 3'h0 == io_c2d_mem_type; // @[Mux.scala 46:19:@3679.4]
  assign mem_type = _T_299 ? 2'h1 : _T_298; // @[Mux.scala 46:16:@3680.4]
  assign _T_301 = 2'h0 == io_c2d_wb_sel; // @[Conditional.scala 37:30:@3685.6]
  assign _T_304 = _T_150 != 5'h0; // @[rvdpath.scala 220:49:@3687.8]
  assign _T_306 = _T_304 ? alu_out : 32'h0; // @[rvdpath.scala 220:40:@3688.8]
  assign _GEN_71 = 5'h0 == _T_150 ? _T_306 : regfile_0; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_72 = 5'h1 == _T_150 ? _T_306 : regfile_1; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_73 = 5'h2 == _T_150 ? _T_306 : regfile_2; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_74 = 5'h3 == _T_150 ? _T_306 : regfile_3; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_75 = 5'h4 == _T_150 ? _T_306 : regfile_4; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_76 = 5'h5 == _T_150 ? _T_306 : regfile_5; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_77 = 5'h6 == _T_150 ? _T_306 : regfile_6; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_78 = 5'h7 == _T_150 ? _T_306 : regfile_7; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_79 = 5'h8 == _T_150 ? _T_306 : regfile_8; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_80 = 5'h9 == _T_150 ? _T_306 : regfile_9; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_81 = 5'ha == _T_150 ? _T_306 : regfile_10; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_82 = 5'hb == _T_150 ? _T_306 : regfile_11; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_83 = 5'hc == _T_150 ? _T_306 : regfile_12; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_84 = 5'hd == _T_150 ? _T_306 : regfile_13; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_85 = 5'he == _T_150 ? _T_306 : regfile_14; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_86 = 5'hf == _T_150 ? _T_306 : regfile_15; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_87 = 5'h10 == _T_150 ? _T_306 : regfile_16; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_88 = 5'h11 == _T_150 ? _T_306 : regfile_17; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_89 = 5'h12 == _T_150 ? _T_306 : regfile_18; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_90 = 5'h13 == _T_150 ? _T_306 : regfile_19; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_91 = 5'h14 == _T_150 ? _T_306 : regfile_20; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_92 = 5'h15 == _T_150 ? _T_306 : regfile_21; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_93 = 5'h16 == _T_150 ? _T_306 : regfile_22; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_94 = 5'h17 == _T_150 ? _T_306 : regfile_23; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_95 = 5'h18 == _T_150 ? _T_306 : regfile_24; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_96 = 5'h19 == _T_150 ? _T_306 : regfile_25; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_97 = 5'h1a == _T_150 ? _T_306 : regfile_26; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_98 = 5'h1b == _T_150 ? _T_306 : regfile_27; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_99 = 5'h1c == _T_150 ? _T_306 : regfile_28; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_100 = 5'h1d == _T_150 ? _T_306 : regfile_29; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_101 = 5'h1e == _T_150 ? _T_306 : regfile_30; // @[rvdpath.scala 220:34:@3689.8]
  assign _GEN_102 = 5'h1f == _T_150 ? _T_306 : regfile_31; // @[rvdpath.scala 220:34:@3689.8]
  assign _T_307 = 2'h1 == io_c2d_wb_sel; // @[Conditional.scala 37:30:@3692.8]
  assign _T_309 = io_dmem_resp_data[7]; // @[rvdpath.scala 228:77:@3695.12]
  assign _T_313 = _T_309 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12:@3697.12]
  assign _T_314 = io_dmem_resp_data[7:0]; // @[rvdpath.scala 228:100:@3698.12]
  assign _T_315 = {_T_313,_T_314}; // @[Cat.scala 30:58:@3699.12]
  assign _T_316 = io_dmem_resp_data[15]; // @[rvdpath.scala 229:77:@3700.12]
  assign _T_320 = _T_316 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@3702.12]
  assign _T_321 = io_dmem_resp_data[15:0]; // @[rvdpath.scala 229:101:@3703.12]
  assign _T_322 = {_T_320,_T_321}; // @[Cat.scala 30:58:@3704.12]
  assign _T_329 = {24'h0,_T_314}; // @[Cat.scala 30:58:@3707.12]
  assign _T_336 = {16'h0,_T_321}; // @[Cat.scala 30:58:@3710.12]
  assign _T_338 = _T_291 ? _T_336 : 32'h0; // @[Mux.scala 46:16:@3712.12]
  assign _T_340 = _T_293 ? _T_329 : _T_338; // @[Mux.scala 46:16:@3714.12]
  assign _T_342 = _T_295 ? io_dmem_resp_data : _T_340; // @[Mux.scala 46:16:@3716.12]
  assign _T_344 = _T_297 ? _T_322 : _T_342; // @[Mux.scala 46:16:@3718.12]
  assign _T_346 = _T_299 ? _T_315 : _T_344; // @[Mux.scala 46:16:@3720.12]
  assign _T_351 = _T_304 ? _T_346 : 32'h0; // @[rvdpath.scala 236:44:@3722.12]
  assign _GEN_103 = 5'h0 == _T_150 ? _T_351 : regfile_0; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_104 = 5'h1 == _T_150 ? _T_351 : regfile_1; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_105 = 5'h2 == _T_150 ? _T_351 : regfile_2; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_106 = 5'h3 == _T_150 ? _T_351 : regfile_3; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_107 = 5'h4 == _T_150 ? _T_351 : regfile_4; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_108 = 5'h5 == _T_150 ? _T_351 : regfile_5; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_109 = 5'h6 == _T_150 ? _T_351 : regfile_6; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_110 = 5'h7 == _T_150 ? _T_351 : regfile_7; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_111 = 5'h8 == _T_150 ? _T_351 : regfile_8; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_112 = 5'h9 == _T_150 ? _T_351 : regfile_9; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_113 = 5'ha == _T_150 ? _T_351 : regfile_10; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_114 = 5'hb == _T_150 ? _T_351 : regfile_11; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_115 = 5'hc == _T_150 ? _T_351 : regfile_12; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_116 = 5'hd == _T_150 ? _T_351 : regfile_13; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_117 = 5'he == _T_150 ? _T_351 : regfile_14; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_118 = 5'hf == _T_150 ? _T_351 : regfile_15; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_119 = 5'h10 == _T_150 ? _T_351 : regfile_16; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_120 = 5'h11 == _T_150 ? _T_351 : regfile_17; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_121 = 5'h12 == _T_150 ? _T_351 : regfile_18; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_122 = 5'h13 == _T_150 ? _T_351 : regfile_19; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_123 = 5'h14 == _T_150 ? _T_351 : regfile_20; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_124 = 5'h15 == _T_150 ? _T_351 : regfile_21; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_125 = 5'h16 == _T_150 ? _T_351 : regfile_22; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_126 = 5'h17 == _T_150 ? _T_351 : regfile_23; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_127 = 5'h18 == _T_150 ? _T_351 : regfile_24; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_128 = 5'h19 == _T_150 ? _T_351 : regfile_25; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_129 = 5'h1a == _T_150 ? _T_351 : regfile_26; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_130 = 5'h1b == _T_150 ? _T_351 : regfile_27; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_131 = 5'h1c == _T_150 ? _T_351 : regfile_28; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_132 = 5'h1d == _T_150 ? _T_351 : regfile_29; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_133 = 5'h1e == _T_150 ? _T_351 : regfile_30; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_134 = 5'h1f == _T_150 ? _T_351 : regfile_31; // @[rvdpath.scala 236:38:@3723.12]
  assign _GEN_135 = io_dmem_resp_valid ? _GEN_103 : regfile_0; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_136 = io_dmem_resp_valid ? _GEN_104 : regfile_1; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_137 = io_dmem_resp_valid ? _GEN_105 : regfile_2; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_138 = io_dmem_resp_valid ? _GEN_106 : regfile_3; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_139 = io_dmem_resp_valid ? _GEN_107 : regfile_4; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_140 = io_dmem_resp_valid ? _GEN_108 : regfile_5; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_141 = io_dmem_resp_valid ? _GEN_109 : regfile_6; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_142 = io_dmem_resp_valid ? _GEN_110 : regfile_7; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_143 = io_dmem_resp_valid ? _GEN_111 : regfile_8; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_144 = io_dmem_resp_valid ? _GEN_112 : regfile_9; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_145 = io_dmem_resp_valid ? _GEN_113 : regfile_10; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_146 = io_dmem_resp_valid ? _GEN_114 : regfile_11; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_147 = io_dmem_resp_valid ? _GEN_115 : regfile_12; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_148 = io_dmem_resp_valid ? _GEN_116 : regfile_13; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_149 = io_dmem_resp_valid ? _GEN_117 : regfile_14; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_150 = io_dmem_resp_valid ? _GEN_118 : regfile_15; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_151 = io_dmem_resp_valid ? _GEN_119 : regfile_16; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_152 = io_dmem_resp_valid ? _GEN_120 : regfile_17; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_153 = io_dmem_resp_valid ? _GEN_121 : regfile_18; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_154 = io_dmem_resp_valid ? _GEN_122 : regfile_19; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_155 = io_dmem_resp_valid ? _GEN_123 : regfile_20; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_156 = io_dmem_resp_valid ? _GEN_124 : regfile_21; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_157 = io_dmem_resp_valid ? _GEN_125 : regfile_22; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_158 = io_dmem_resp_valid ? _GEN_126 : regfile_23; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_159 = io_dmem_resp_valid ? _GEN_127 : regfile_24; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_160 = io_dmem_resp_valid ? _GEN_128 : regfile_25; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_161 = io_dmem_resp_valid ? _GEN_129 : regfile_26; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_162 = io_dmem_resp_valid ? _GEN_130 : regfile_27; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_163 = io_dmem_resp_valid ? _GEN_131 : regfile_28; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_164 = io_dmem_resp_valid ? _GEN_132 : regfile_29; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_165 = io_dmem_resp_valid ? _GEN_133 : regfile_30; // @[rvdpath.scala 223:42:@3694.10]
  assign _GEN_166 = io_dmem_resp_valid ? _GEN_134 : regfile_31; // @[rvdpath.scala 223:42:@3694.10]
  assign _T_352 = 2'h2 == io_c2d_wb_sel; // @[Conditional.scala 37:30:@3727.10]
  assign _T_357 = _T_304 ? pc_a4 : 32'h0; // @[rvdpath.scala 241:40:@3730.12]
  assign _GEN_167 = 5'h0 == _T_150 ? _T_357 : regfile_0; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_168 = 5'h1 == _T_150 ? _T_357 : regfile_1; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_169 = 5'h2 == _T_150 ? _T_357 : regfile_2; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_170 = 5'h3 == _T_150 ? _T_357 : regfile_3; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_171 = 5'h4 == _T_150 ? _T_357 : regfile_4; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_172 = 5'h5 == _T_150 ? _T_357 : regfile_5; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_173 = 5'h6 == _T_150 ? _T_357 : regfile_6; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_174 = 5'h7 == _T_150 ? _T_357 : regfile_7; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_175 = 5'h8 == _T_150 ? _T_357 : regfile_8; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_176 = 5'h9 == _T_150 ? _T_357 : regfile_9; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_177 = 5'ha == _T_150 ? _T_357 : regfile_10; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_178 = 5'hb == _T_150 ? _T_357 : regfile_11; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_179 = 5'hc == _T_150 ? _T_357 : regfile_12; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_180 = 5'hd == _T_150 ? _T_357 : regfile_13; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_181 = 5'he == _T_150 ? _T_357 : regfile_14; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_182 = 5'hf == _T_150 ? _T_357 : regfile_15; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_183 = 5'h10 == _T_150 ? _T_357 : regfile_16; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_184 = 5'h11 == _T_150 ? _T_357 : regfile_17; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_185 = 5'h12 == _T_150 ? _T_357 : regfile_18; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_186 = 5'h13 == _T_150 ? _T_357 : regfile_19; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_187 = 5'h14 == _T_150 ? _T_357 : regfile_20; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_188 = 5'h15 == _T_150 ? _T_357 : regfile_21; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_189 = 5'h16 == _T_150 ? _T_357 : regfile_22; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_190 = 5'h17 == _T_150 ? _T_357 : regfile_23; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_191 = 5'h18 == _T_150 ? _T_357 : regfile_24; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_192 = 5'h19 == _T_150 ? _T_357 : regfile_25; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_193 = 5'h1a == _T_150 ? _T_357 : regfile_26; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_194 = 5'h1b == _T_150 ? _T_357 : regfile_27; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_195 = 5'h1c == _T_150 ? _T_357 : regfile_28; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_196 = 5'h1d == _T_150 ? _T_357 : regfile_29; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_197 = 5'h1e == _T_150 ? _T_357 : regfile_30; // @[rvdpath.scala 241:34:@3731.12]
  assign _GEN_198 = 5'h1f == _T_150 ? _T_357 : regfile_31; // @[rvdpath.scala 241:34:@3731.12]
  assign _T_358 = 2'h3 == io_c2d_wb_sel; // @[Conditional.scala 37:30:@3734.12]
  assign csr_rdata = csr_io_rdata; // @[rvdpath.scala 192:25:@3664.4]
  assign _T_363 = _T_304 ? csr_rdata : 32'h0; // @[rvdpath.scala 245:40:@3737.14]
  assign _GEN_199 = 5'h0 == _T_150 ? _T_363 : regfile_0; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_200 = 5'h1 == _T_150 ? _T_363 : regfile_1; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_201 = 5'h2 == _T_150 ? _T_363 : regfile_2; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_202 = 5'h3 == _T_150 ? _T_363 : regfile_3; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_203 = 5'h4 == _T_150 ? _T_363 : regfile_4; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_204 = 5'h5 == _T_150 ? _T_363 : regfile_5; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_205 = 5'h6 == _T_150 ? _T_363 : regfile_6; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_206 = 5'h7 == _T_150 ? _T_363 : regfile_7; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_207 = 5'h8 == _T_150 ? _T_363 : regfile_8; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_208 = 5'h9 == _T_150 ? _T_363 : regfile_9; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_209 = 5'ha == _T_150 ? _T_363 : regfile_10; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_210 = 5'hb == _T_150 ? _T_363 : regfile_11; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_211 = 5'hc == _T_150 ? _T_363 : regfile_12; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_212 = 5'hd == _T_150 ? _T_363 : regfile_13; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_213 = 5'he == _T_150 ? _T_363 : regfile_14; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_214 = 5'hf == _T_150 ? _T_363 : regfile_15; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_215 = 5'h10 == _T_150 ? _T_363 : regfile_16; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_216 = 5'h11 == _T_150 ? _T_363 : regfile_17; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_217 = 5'h12 == _T_150 ? _T_363 : regfile_18; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_218 = 5'h13 == _T_150 ? _T_363 : regfile_19; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_219 = 5'h14 == _T_150 ? _T_363 : regfile_20; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_220 = 5'h15 == _T_150 ? _T_363 : regfile_21; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_221 = 5'h16 == _T_150 ? _T_363 : regfile_22; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_222 = 5'h17 == _T_150 ? _T_363 : regfile_23; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_223 = 5'h18 == _T_150 ? _T_363 : regfile_24; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_224 = 5'h19 == _T_150 ? _T_363 : regfile_25; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_225 = 5'h1a == _T_150 ? _T_363 : regfile_26; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_226 = 5'h1b == _T_150 ? _T_363 : regfile_27; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_227 = 5'h1c == _T_150 ? _T_363 : regfile_28; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_228 = 5'h1d == _T_150 ? _T_363 : regfile_29; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_229 = 5'h1e == _T_150 ? _T_363 : regfile_30; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_230 = 5'h1f == _T_150 ? _T_363 : regfile_31; // @[rvdpath.scala 245:34:@3738.14]
  assign _GEN_231 = _T_358 ? _GEN_199 : regfile_0; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_232 = _T_358 ? _GEN_200 : regfile_1; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_233 = _T_358 ? _GEN_201 : regfile_2; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_234 = _T_358 ? _GEN_202 : regfile_3; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_235 = _T_358 ? _GEN_203 : regfile_4; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_236 = _T_358 ? _GEN_204 : regfile_5; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_237 = _T_358 ? _GEN_205 : regfile_6; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_238 = _T_358 ? _GEN_206 : regfile_7; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_239 = _T_358 ? _GEN_207 : regfile_8; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_240 = _T_358 ? _GEN_208 : regfile_9; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_241 = _T_358 ? _GEN_209 : regfile_10; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_242 = _T_358 ? _GEN_210 : regfile_11; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_243 = _T_358 ? _GEN_211 : regfile_12; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_244 = _T_358 ? _GEN_212 : regfile_13; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_245 = _T_358 ? _GEN_213 : regfile_14; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_246 = _T_358 ? _GEN_214 : regfile_15; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_247 = _T_358 ? _GEN_215 : regfile_16; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_248 = _T_358 ? _GEN_216 : regfile_17; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_249 = _T_358 ? _GEN_217 : regfile_18; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_250 = _T_358 ? _GEN_218 : regfile_19; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_251 = _T_358 ? _GEN_219 : regfile_20; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_252 = _T_358 ? _GEN_220 : regfile_21; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_253 = _T_358 ? _GEN_221 : regfile_22; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_254 = _T_358 ? _GEN_222 : regfile_23; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_255 = _T_358 ? _GEN_223 : regfile_24; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_256 = _T_358 ? _GEN_224 : regfile_25; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_257 = _T_358 ? _GEN_225 : regfile_26; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_258 = _T_358 ? _GEN_226 : regfile_27; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_259 = _T_358 ? _GEN_227 : regfile_28; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_260 = _T_358 ? _GEN_228 : regfile_29; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_261 = _T_358 ? _GEN_229 : regfile_30; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_262 = _T_358 ? _GEN_230 : regfile_31; // @[Conditional.scala 39:67:@3735.12]
  assign _GEN_263 = _T_352 ? _GEN_167 : _GEN_231; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_264 = _T_352 ? _GEN_168 : _GEN_232; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_265 = _T_352 ? _GEN_169 : _GEN_233; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_266 = _T_352 ? _GEN_170 : _GEN_234; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_267 = _T_352 ? _GEN_171 : _GEN_235; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_268 = _T_352 ? _GEN_172 : _GEN_236; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_269 = _T_352 ? _GEN_173 : _GEN_237; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_270 = _T_352 ? _GEN_174 : _GEN_238; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_271 = _T_352 ? _GEN_175 : _GEN_239; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_272 = _T_352 ? _GEN_176 : _GEN_240; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_273 = _T_352 ? _GEN_177 : _GEN_241; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_274 = _T_352 ? _GEN_178 : _GEN_242; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_275 = _T_352 ? _GEN_179 : _GEN_243; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_276 = _T_352 ? _GEN_180 : _GEN_244; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_277 = _T_352 ? _GEN_181 : _GEN_245; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_278 = _T_352 ? _GEN_182 : _GEN_246; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_279 = _T_352 ? _GEN_183 : _GEN_247; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_280 = _T_352 ? _GEN_184 : _GEN_248; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_281 = _T_352 ? _GEN_185 : _GEN_249; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_282 = _T_352 ? _GEN_186 : _GEN_250; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_283 = _T_352 ? _GEN_187 : _GEN_251; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_284 = _T_352 ? _GEN_188 : _GEN_252; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_285 = _T_352 ? _GEN_189 : _GEN_253; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_286 = _T_352 ? _GEN_190 : _GEN_254; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_287 = _T_352 ? _GEN_191 : _GEN_255; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_288 = _T_352 ? _GEN_192 : _GEN_256; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_289 = _T_352 ? _GEN_193 : _GEN_257; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_290 = _T_352 ? _GEN_194 : _GEN_258; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_291 = _T_352 ? _GEN_195 : _GEN_259; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_292 = _T_352 ? _GEN_196 : _GEN_260; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_293 = _T_352 ? _GEN_197 : _GEN_261; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_294 = _T_352 ? _GEN_198 : _GEN_262; // @[Conditional.scala 39:67:@3728.10]
  assign _GEN_295 = _T_307 ? _GEN_135 : _GEN_263; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_296 = _T_307 ? _GEN_136 : _GEN_264; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_297 = _T_307 ? _GEN_137 : _GEN_265; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_298 = _T_307 ? _GEN_138 : _GEN_266; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_299 = _T_307 ? _GEN_139 : _GEN_267; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_300 = _T_307 ? _GEN_140 : _GEN_268; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_301 = _T_307 ? _GEN_141 : _GEN_269; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_302 = _T_307 ? _GEN_142 : _GEN_270; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_303 = _T_307 ? _GEN_143 : _GEN_271; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_304 = _T_307 ? _GEN_144 : _GEN_272; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_305 = _T_307 ? _GEN_145 : _GEN_273; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_306 = _T_307 ? _GEN_146 : _GEN_274; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_307 = _T_307 ? _GEN_147 : _GEN_275; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_308 = _T_307 ? _GEN_148 : _GEN_276; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_309 = _T_307 ? _GEN_149 : _GEN_277; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_310 = _T_307 ? _GEN_150 : _GEN_278; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_311 = _T_307 ? _GEN_151 : _GEN_279; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_312 = _T_307 ? _GEN_152 : _GEN_280; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_313 = _T_307 ? _GEN_153 : _GEN_281; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_314 = _T_307 ? _GEN_154 : _GEN_282; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_315 = _T_307 ? _GEN_155 : _GEN_283; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_316 = _T_307 ? _GEN_156 : _GEN_284; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_317 = _T_307 ? _GEN_157 : _GEN_285; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_318 = _T_307 ? _GEN_158 : _GEN_286; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_319 = _T_307 ? _GEN_159 : _GEN_287; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_320 = _T_307 ? _GEN_160 : _GEN_288; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_321 = _T_307 ? _GEN_161 : _GEN_289; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_322 = _T_307 ? _GEN_162 : _GEN_290; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_323 = _T_307 ? _GEN_163 : _GEN_291; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_324 = _T_307 ? _GEN_164 : _GEN_292; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_325 = _T_307 ? _GEN_165 : _GEN_293; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_326 = _T_307 ? _GEN_166 : _GEN_294; // @[Conditional.scala 39:67:@3693.8]
  assign _GEN_327 = _T_301 ? _GEN_71 : _GEN_295; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_328 = _T_301 ? _GEN_72 : _GEN_296; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_329 = _T_301 ? _GEN_73 : _GEN_297; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_330 = _T_301 ? _GEN_74 : _GEN_298; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_331 = _T_301 ? _GEN_75 : _GEN_299; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_332 = _T_301 ? _GEN_76 : _GEN_300; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_333 = _T_301 ? _GEN_77 : _GEN_301; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_334 = _T_301 ? _GEN_78 : _GEN_302; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_335 = _T_301 ? _GEN_79 : _GEN_303; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_336 = _T_301 ? _GEN_80 : _GEN_304; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_337 = _T_301 ? _GEN_81 : _GEN_305; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_338 = _T_301 ? _GEN_82 : _GEN_306; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_339 = _T_301 ? _GEN_83 : _GEN_307; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_340 = _T_301 ? _GEN_84 : _GEN_308; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_341 = _T_301 ? _GEN_85 : _GEN_309; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_342 = _T_301 ? _GEN_86 : _GEN_310; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_343 = _T_301 ? _GEN_87 : _GEN_311; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_344 = _T_301 ? _GEN_88 : _GEN_312; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_345 = _T_301 ? _GEN_89 : _GEN_313; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_346 = _T_301 ? _GEN_90 : _GEN_314; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_347 = _T_301 ? _GEN_91 : _GEN_315; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_348 = _T_301 ? _GEN_92 : _GEN_316; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_349 = _T_301 ? _GEN_93 : _GEN_317; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_350 = _T_301 ? _GEN_94 : _GEN_318; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_351 = _T_301 ? _GEN_95 : _GEN_319; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_352 = _T_301 ? _GEN_96 : _GEN_320; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_353 = _T_301 ? _GEN_97 : _GEN_321; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_354 = _T_301 ? _GEN_98 : _GEN_322; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_355 = _T_301 ? _GEN_99 : _GEN_323; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_356 = _T_301 ? _GEN_100 : _GEN_324; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_357 = _T_301 ? _GEN_101 : _GEN_325; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_358 = _T_301 ? _GEN_102 : _GEN_326; // @[Conditional.scala 40:58:@3686.6]
  assign _GEN_359 = io_c2d_reg_wren ? _GEN_327 : regfile_0; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_360 = io_c2d_reg_wren ? _GEN_328 : regfile_1; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_361 = io_c2d_reg_wren ? _GEN_329 : regfile_2; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_362 = io_c2d_reg_wren ? _GEN_330 : regfile_3; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_363 = io_c2d_reg_wren ? _GEN_331 : regfile_4; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_364 = io_c2d_reg_wren ? _GEN_332 : regfile_5; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_365 = io_c2d_reg_wren ? _GEN_333 : regfile_6; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_366 = io_c2d_reg_wren ? _GEN_334 : regfile_7; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_367 = io_c2d_reg_wren ? _GEN_335 : regfile_8; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_368 = io_c2d_reg_wren ? _GEN_336 : regfile_9; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_369 = io_c2d_reg_wren ? _GEN_337 : regfile_10; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_370 = io_c2d_reg_wren ? _GEN_338 : regfile_11; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_371 = io_c2d_reg_wren ? _GEN_339 : regfile_12; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_372 = io_c2d_reg_wren ? _GEN_340 : regfile_13; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_373 = io_c2d_reg_wren ? _GEN_341 : regfile_14; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_374 = io_c2d_reg_wren ? _GEN_342 : regfile_15; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_375 = io_c2d_reg_wren ? _GEN_343 : regfile_16; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_376 = io_c2d_reg_wren ? _GEN_344 : regfile_17; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_377 = io_c2d_reg_wren ? _GEN_345 : regfile_18; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_378 = io_c2d_reg_wren ? _GEN_346 : regfile_19; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_379 = io_c2d_reg_wren ? _GEN_347 : regfile_20; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_380 = io_c2d_reg_wren ? _GEN_348 : regfile_21; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_381 = io_c2d_reg_wren ? _GEN_349 : regfile_22; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_382 = io_c2d_reg_wren ? _GEN_350 : regfile_23; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_383 = io_c2d_reg_wren ? _GEN_351 : regfile_24; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_384 = io_c2d_reg_wren ? _GEN_352 : regfile_25; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_385 = io_c2d_reg_wren ? _GEN_353 : regfile_26; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_386 = io_c2d_reg_wren ? _GEN_354 : regfile_27; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_387 = io_c2d_reg_wren ? _GEN_355 : regfile_28; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_388 = io_c2d_reg_wren ? _GEN_356 : regfile_29; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_389 = io_c2d_reg_wren ? _GEN_357 : regfile_30; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_390 = io_c2d_reg_wren ? _GEN_358 : regfile_31; // @[rvdpath.scala 216:47:@3684.4]
  assign _GEN_391 = 5'h1 == io_ddpath_addr ? regfile_1 : regfile_0; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_392 = 5'h2 == io_ddpath_addr ? regfile_2 : _GEN_391; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_393 = 5'h3 == io_ddpath_addr ? regfile_3 : _GEN_392; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_394 = 5'h4 == io_ddpath_addr ? regfile_4 : _GEN_393; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_395 = 5'h5 == io_ddpath_addr ? regfile_5 : _GEN_394; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_396 = 5'h6 == io_ddpath_addr ? regfile_6 : _GEN_395; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_397 = 5'h7 == io_ddpath_addr ? regfile_7 : _GEN_396; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_398 = 5'h8 == io_ddpath_addr ? regfile_8 : _GEN_397; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_399 = 5'h9 == io_ddpath_addr ? regfile_9 : _GEN_398; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_400 = 5'ha == io_ddpath_addr ? regfile_10 : _GEN_399; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_401 = 5'hb == io_ddpath_addr ? regfile_11 : _GEN_400; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_402 = 5'hc == io_ddpath_addr ? regfile_12 : _GEN_401; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_403 = 5'hd == io_ddpath_addr ? regfile_13 : _GEN_402; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_404 = 5'he == io_ddpath_addr ? regfile_14 : _GEN_403; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_405 = 5'hf == io_ddpath_addr ? regfile_15 : _GEN_404; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_406 = 5'h10 == io_ddpath_addr ? regfile_16 : _GEN_405; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_407 = 5'h11 == io_ddpath_addr ? regfile_17 : _GEN_406; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_408 = 5'h12 == io_ddpath_addr ? regfile_18 : _GEN_407; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_409 = 5'h13 == io_ddpath_addr ? regfile_19 : _GEN_408; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_410 = 5'h14 == io_ddpath_addr ? regfile_20 : _GEN_409; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_411 = 5'h15 == io_ddpath_addr ? regfile_21 : _GEN_410; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_412 = 5'h16 == io_ddpath_addr ? regfile_22 : _GEN_411; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_413 = 5'h17 == io_ddpath_addr ? regfile_23 : _GEN_412; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_414 = 5'h18 == io_ddpath_addr ? regfile_24 : _GEN_413; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_415 = 5'h19 == io_ddpath_addr ? regfile_25 : _GEN_414; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_416 = 5'h1a == io_ddpath_addr ? regfile_26 : _GEN_415; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_417 = 5'h1b == io_ddpath_addr ? regfile_27 : _GEN_416; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_418 = 5'h1c == io_ddpath_addr ? regfile_28 : _GEN_417; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_419 = 5'h1d == io_ddpath_addr ? regfile_29 : _GEN_418; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_420 = 5'h1e == io_ddpath_addr ? regfile_30 : _GEN_419; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_421 = 5'h1f == io_ddpath_addr ? regfile_31 : _GEN_420; // @[rvdpath.scala 265:21:@3755.4]
  assign _GEN_422 = 5'h0 == io_ddpath_addr ? io_ddpath_wdata : _GEN_359; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_423 = 5'h1 == io_ddpath_addr ? io_ddpath_wdata : _GEN_360; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_424 = 5'h2 == io_ddpath_addr ? io_ddpath_wdata : _GEN_361; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_425 = 5'h3 == io_ddpath_addr ? io_ddpath_wdata : _GEN_362; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_426 = 5'h4 == io_ddpath_addr ? io_ddpath_wdata : _GEN_363; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_427 = 5'h5 == io_ddpath_addr ? io_ddpath_wdata : _GEN_364; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_428 = 5'h6 == io_ddpath_addr ? io_ddpath_wdata : _GEN_365; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_429 = 5'h7 == io_ddpath_addr ? io_ddpath_wdata : _GEN_366; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_430 = 5'h8 == io_ddpath_addr ? io_ddpath_wdata : _GEN_367; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_431 = 5'h9 == io_ddpath_addr ? io_ddpath_wdata : _GEN_368; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_432 = 5'ha == io_ddpath_addr ? io_ddpath_wdata : _GEN_369; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_433 = 5'hb == io_ddpath_addr ? io_ddpath_wdata : _GEN_370; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_434 = 5'hc == io_ddpath_addr ? io_ddpath_wdata : _GEN_371; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_435 = 5'hd == io_ddpath_addr ? io_ddpath_wdata : _GEN_372; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_436 = 5'he == io_ddpath_addr ? io_ddpath_wdata : _GEN_373; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_437 = 5'hf == io_ddpath_addr ? io_ddpath_wdata : _GEN_374; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_438 = 5'h10 == io_ddpath_addr ? io_ddpath_wdata : _GEN_375; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_439 = 5'h11 == io_ddpath_addr ? io_ddpath_wdata : _GEN_376; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_440 = 5'h12 == io_ddpath_addr ? io_ddpath_wdata : _GEN_377; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_441 = 5'h13 == io_ddpath_addr ? io_ddpath_wdata : _GEN_378; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_442 = 5'h14 == io_ddpath_addr ? io_ddpath_wdata : _GEN_379; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_443 = 5'h15 == io_ddpath_addr ? io_ddpath_wdata : _GEN_380; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_444 = 5'h16 == io_ddpath_addr ? io_ddpath_wdata : _GEN_381; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_445 = 5'h17 == io_ddpath_addr ? io_ddpath_wdata : _GEN_382; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_446 = 5'h18 == io_ddpath_addr ? io_ddpath_wdata : _GEN_383; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_447 = 5'h19 == io_ddpath_addr ? io_ddpath_wdata : _GEN_384; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_448 = 5'h1a == io_ddpath_addr ? io_ddpath_wdata : _GEN_385; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_449 = 5'h1b == io_ddpath_addr ? io_ddpath_wdata : _GEN_386; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_450 = 5'h1c == io_ddpath_addr ? io_ddpath_wdata : _GEN_387; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_451 = 5'h1d == io_ddpath_addr ? io_ddpath_wdata : _GEN_388; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_452 = 5'h1e == io_ddpath_addr ? io_ddpath_wdata : _GEN_389; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_453 = 5'h1f == io_ddpath_addr ? io_ddpath_wdata : _GEN_390; // @[rvdpath.scala 267:33:@3757.6]
  assign _GEN_454 = io_ddpath_valid ? _GEN_422 : _GEN_359; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_455 = io_ddpath_valid ? _GEN_423 : _GEN_360; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_456 = io_ddpath_valid ? _GEN_424 : _GEN_361; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_457 = io_ddpath_valid ? _GEN_425 : _GEN_362; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_458 = io_ddpath_valid ? _GEN_426 : _GEN_363; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_459 = io_ddpath_valid ? _GEN_427 : _GEN_364; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_460 = io_ddpath_valid ? _GEN_428 : _GEN_365; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_461 = io_ddpath_valid ? _GEN_429 : _GEN_366; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_462 = io_ddpath_valid ? _GEN_430 : _GEN_367; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_463 = io_ddpath_valid ? _GEN_431 : _GEN_368; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_464 = io_ddpath_valid ? _GEN_432 : _GEN_369; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_465 = io_ddpath_valid ? _GEN_433 : _GEN_370; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_466 = io_ddpath_valid ? _GEN_434 : _GEN_371; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_467 = io_ddpath_valid ? _GEN_435 : _GEN_372; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_468 = io_ddpath_valid ? _GEN_436 : _GEN_373; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_469 = io_ddpath_valid ? _GEN_437 : _GEN_374; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_470 = io_ddpath_valid ? _GEN_438 : _GEN_375; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_471 = io_ddpath_valid ? _GEN_439 : _GEN_376; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_472 = io_ddpath_valid ? _GEN_440 : _GEN_377; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_473 = io_ddpath_valid ? _GEN_441 : _GEN_378; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_474 = io_ddpath_valid ? _GEN_442 : _GEN_379; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_475 = io_ddpath_valid ? _GEN_443 : _GEN_380; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_476 = io_ddpath_valid ? _GEN_444 : _GEN_381; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_477 = io_ddpath_valid ? _GEN_445 : _GEN_382; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_478 = io_ddpath_valid ? _GEN_446 : _GEN_383; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_479 = io_ddpath_valid ? _GEN_447 : _GEN_384; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_480 = io_ddpath_valid ? _GEN_448 : _GEN_385; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_481 = io_ddpath_valid ? _GEN_449 : _GEN_386; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_482 = io_ddpath_valid ? _GEN_450 : _GEN_387; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_483 = io_ddpath_valid ? _GEN_451 : _GEN_388; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_484 = io_ddpath_valid ? _GEN_452 : _GEN_389; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_485 = io_ddpath_valid ? _GEN_453 : _GEN_390; // @[rvdpath.scala 266:26:@3756.4]
  assign _GEN_486 = reset ? 32'h80000000 : _GEN_8; // @[rvdpath.scala 271:26:@3760.4]
  assign _GEN_487 = reset ? 1'h0 : 1'h1; // @[rvdpath.scala 271:26:@3760.4]
  assign _GEN_488 = reset ? 1'h0 : io_c2d_mem_en; // @[rvdpath.scala 271:26:@3760.4]
  assign io_imem_req_addr = pc;
  assign io_imem_req_valid = _GEN_487;
  assign io_dmem_req_addr = alu_out;
  assign io_dmem_req_data = rs2_data;
  assign io_dmem_req_mfunc = io_c2d_mem_wren;
  assign io_dmem_req_mtype = mem_type;
  assign io_dmem_req_valid = _GEN_488;
  assign io_d2c_inst = inst;
  assign io_d2c_dexcp = csr_io_csr_excp;
  assign io_ddpath_rdata = _GEN_421;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_addr = _T_143;
  assign csr_io_wdata = alu_opd1;
  assign csr_io_op = io_c2d_csr_cmd;
  assign csr_io_core_pc = pc;
  assign csr_io_core_excp = io_c2d_cexcp;
  assign csr_io_core_cause = io_c2d_ccause;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  regfile_0 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  regfile_1 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  regfile_2 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  regfile_3 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  regfile_4 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  regfile_5 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  regfile_6 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  regfile_7 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  regfile_8 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  regfile_9 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  regfile_10 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  regfile_11 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  regfile_12 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  regfile_13 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  regfile_14 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  regfile_15 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  regfile_16 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  regfile_17 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  regfile_18 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  regfile_19 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  regfile_20 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  regfile_21 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  regfile_22 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  regfile_23 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  regfile_24 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  regfile_25 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  regfile_26 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  regfile_27 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  regfile_28 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  regfile_29 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  regfile_30 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  regfile_31 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h80000000;
    end else begin
      if (pc_update) begin
        if (_T_79) begin
          pc <= pc_a4;
        end else begin
          if (_T_77) begin
            if (_T_285) begin
              if (bcmp_eq) begin
                pc <= alu_out;
              end else begin
                pc <= pc_a4;
              end
            end else begin
              if (_T_283) begin
                if (_T_265) begin
                  pc <= alu_out;
                end else begin
                  pc <= pc_a4;
                end
              end else begin
                if (_T_281) begin
                  if (bcmp_lt) begin
                    pc <= alu_out;
                  end else begin
                    pc <= pc_a4;
                  end
                end else begin
                  if (_T_279) begin
                    if (_T_269) begin
                      pc <= alu_out;
                    end else begin
                      pc <= pc_a4;
                    end
                  end else begin
                    if (_T_277) begin
                      if (bcmp_ltu) begin
                        pc <= alu_out;
                      end else begin
                        pc <= pc_a4;
                      end
                    end else begin
                      if (_T_275) begin
                        if (_T_273) begin
                          pc <= alu_out;
                        end else begin
                          pc <= pc_a4;
                        end
                      end else begin
                        pc <= pc_a4;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_75) begin
              pc <= alu_out;
            end else begin
              if (_T_73) begin
                pc <= pc_ex;
              end else begin
                pc <= pc_a4;
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h0 == io_ddpath_addr) begin
        regfile_0 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h0 == _T_150) begin
              if (_T_304) begin
                regfile_0 <= alu_out;
              end else begin
                regfile_0 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h0 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_0 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_0 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_0 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_0 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_0 <= _T_336;
                            end else begin
                              regfile_0 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_0 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h0 == _T_150) begin
                  if (_T_304) begin
                    regfile_0 <= pc_a4;
                  end else begin
                    regfile_0 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h0 == _T_150) begin
                    if (_T_304) begin
                      regfile_0 <= csr_rdata;
                    end else begin
                      regfile_0 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h0 == _T_150) begin
            if (_T_304) begin
              regfile_0 <= alu_out;
            end else begin
              regfile_0 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h0 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_0 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_0 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_0 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_0 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_0 <= _T_336;
                          end else begin
                            regfile_0 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_0 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h0 == _T_150) begin
                if (_T_304) begin
                  regfile_0 <= pc_a4;
                end else begin
                  regfile_0 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h0 == _T_150) begin
                  if (_T_304) begin
                    regfile_0 <= csr_rdata;
                  end else begin
                    regfile_0 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h1 == io_ddpath_addr) begin
        regfile_1 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h1 == _T_150) begin
              if (_T_304) begin
                regfile_1 <= alu_out;
              end else begin
                regfile_1 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h1 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_1 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_1 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_1 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_1 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_1 <= _T_336;
                            end else begin
                              regfile_1 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_1 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h1 == _T_150) begin
                  if (_T_304) begin
                    regfile_1 <= pc_a4;
                  end else begin
                    regfile_1 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h1 == _T_150) begin
                    if (_T_304) begin
                      regfile_1 <= csr_rdata;
                    end else begin
                      regfile_1 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h1 == _T_150) begin
            if (_T_304) begin
              regfile_1 <= alu_out;
            end else begin
              regfile_1 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h1 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_1 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_1 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_1 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_1 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_1 <= _T_336;
                          end else begin
                            regfile_1 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_1 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h1 == _T_150) begin
                if (_T_304) begin
                  regfile_1 <= pc_a4;
                end else begin
                  regfile_1 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h1 == _T_150) begin
                  if (_T_304) begin
                    regfile_1 <= csr_rdata;
                  end else begin
                    regfile_1 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h2 == io_ddpath_addr) begin
        regfile_2 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h2 == _T_150) begin
              if (_T_304) begin
                regfile_2 <= alu_out;
              end else begin
                regfile_2 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h2 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_2 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_2 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_2 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_2 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_2 <= _T_336;
                            end else begin
                              regfile_2 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_2 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h2 == _T_150) begin
                  if (_T_304) begin
                    regfile_2 <= pc_a4;
                  end else begin
                    regfile_2 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h2 == _T_150) begin
                    if (_T_304) begin
                      regfile_2 <= csr_rdata;
                    end else begin
                      regfile_2 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h2 == _T_150) begin
            if (_T_304) begin
              regfile_2 <= alu_out;
            end else begin
              regfile_2 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h2 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_2 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_2 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_2 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_2 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_2 <= _T_336;
                          end else begin
                            regfile_2 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_2 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h2 == _T_150) begin
                if (_T_304) begin
                  regfile_2 <= pc_a4;
                end else begin
                  regfile_2 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h2 == _T_150) begin
                  if (_T_304) begin
                    regfile_2 <= csr_rdata;
                  end else begin
                    regfile_2 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h3 == io_ddpath_addr) begin
        regfile_3 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h3 == _T_150) begin
              if (_T_304) begin
                regfile_3 <= alu_out;
              end else begin
                regfile_3 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h3 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_3 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_3 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_3 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_3 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_3 <= _T_336;
                            end else begin
                              regfile_3 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_3 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h3 == _T_150) begin
                  if (_T_304) begin
                    regfile_3 <= pc_a4;
                  end else begin
                    regfile_3 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h3 == _T_150) begin
                    if (_T_304) begin
                      regfile_3 <= csr_rdata;
                    end else begin
                      regfile_3 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h3 == _T_150) begin
            if (_T_304) begin
              regfile_3 <= alu_out;
            end else begin
              regfile_3 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h3 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_3 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_3 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_3 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_3 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_3 <= _T_336;
                          end else begin
                            regfile_3 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_3 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h3 == _T_150) begin
                if (_T_304) begin
                  regfile_3 <= pc_a4;
                end else begin
                  regfile_3 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h3 == _T_150) begin
                  if (_T_304) begin
                    regfile_3 <= csr_rdata;
                  end else begin
                    regfile_3 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h4 == io_ddpath_addr) begin
        regfile_4 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h4 == _T_150) begin
              if (_T_304) begin
                regfile_4 <= alu_out;
              end else begin
                regfile_4 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h4 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_4 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_4 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_4 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_4 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_4 <= _T_336;
                            end else begin
                              regfile_4 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_4 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h4 == _T_150) begin
                  if (_T_304) begin
                    regfile_4 <= pc_a4;
                  end else begin
                    regfile_4 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h4 == _T_150) begin
                    if (_T_304) begin
                      regfile_4 <= csr_rdata;
                    end else begin
                      regfile_4 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h4 == _T_150) begin
            if (_T_304) begin
              regfile_4 <= alu_out;
            end else begin
              regfile_4 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h4 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_4 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_4 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_4 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_4 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_4 <= _T_336;
                          end else begin
                            regfile_4 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_4 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h4 == _T_150) begin
                if (_T_304) begin
                  regfile_4 <= pc_a4;
                end else begin
                  regfile_4 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h4 == _T_150) begin
                  if (_T_304) begin
                    regfile_4 <= csr_rdata;
                  end else begin
                    regfile_4 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h5 == io_ddpath_addr) begin
        regfile_5 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h5 == _T_150) begin
              if (_T_304) begin
                regfile_5 <= alu_out;
              end else begin
                regfile_5 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h5 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_5 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_5 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_5 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_5 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_5 <= _T_336;
                            end else begin
                              regfile_5 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_5 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h5 == _T_150) begin
                  if (_T_304) begin
                    regfile_5 <= pc_a4;
                  end else begin
                    regfile_5 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h5 == _T_150) begin
                    if (_T_304) begin
                      regfile_5 <= csr_rdata;
                    end else begin
                      regfile_5 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h5 == _T_150) begin
            if (_T_304) begin
              regfile_5 <= alu_out;
            end else begin
              regfile_5 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h5 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_5 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_5 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_5 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_5 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_5 <= _T_336;
                          end else begin
                            regfile_5 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_5 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h5 == _T_150) begin
                if (_T_304) begin
                  regfile_5 <= pc_a4;
                end else begin
                  regfile_5 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h5 == _T_150) begin
                  if (_T_304) begin
                    regfile_5 <= csr_rdata;
                  end else begin
                    regfile_5 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h6 == io_ddpath_addr) begin
        regfile_6 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h6 == _T_150) begin
              if (_T_304) begin
                regfile_6 <= alu_out;
              end else begin
                regfile_6 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h6 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_6 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_6 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_6 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_6 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_6 <= _T_336;
                            end else begin
                              regfile_6 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_6 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h6 == _T_150) begin
                  if (_T_304) begin
                    regfile_6 <= pc_a4;
                  end else begin
                    regfile_6 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h6 == _T_150) begin
                    if (_T_304) begin
                      regfile_6 <= csr_rdata;
                    end else begin
                      regfile_6 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h6 == _T_150) begin
            if (_T_304) begin
              regfile_6 <= alu_out;
            end else begin
              regfile_6 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h6 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_6 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_6 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_6 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_6 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_6 <= _T_336;
                          end else begin
                            regfile_6 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_6 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h6 == _T_150) begin
                if (_T_304) begin
                  regfile_6 <= pc_a4;
                end else begin
                  regfile_6 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h6 == _T_150) begin
                  if (_T_304) begin
                    regfile_6 <= csr_rdata;
                  end else begin
                    regfile_6 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h7 == io_ddpath_addr) begin
        regfile_7 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h7 == _T_150) begin
              if (_T_304) begin
                regfile_7 <= alu_out;
              end else begin
                regfile_7 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h7 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_7 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_7 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_7 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_7 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_7 <= _T_336;
                            end else begin
                              regfile_7 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_7 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h7 == _T_150) begin
                  if (_T_304) begin
                    regfile_7 <= pc_a4;
                  end else begin
                    regfile_7 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h7 == _T_150) begin
                    if (_T_304) begin
                      regfile_7 <= csr_rdata;
                    end else begin
                      regfile_7 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h7 == _T_150) begin
            if (_T_304) begin
              regfile_7 <= alu_out;
            end else begin
              regfile_7 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h7 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_7 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_7 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_7 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_7 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_7 <= _T_336;
                          end else begin
                            regfile_7 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_7 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h7 == _T_150) begin
                if (_T_304) begin
                  regfile_7 <= pc_a4;
                end else begin
                  regfile_7 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h7 == _T_150) begin
                  if (_T_304) begin
                    regfile_7 <= csr_rdata;
                  end else begin
                    regfile_7 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h8 == io_ddpath_addr) begin
        regfile_8 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h8 == _T_150) begin
              if (_T_304) begin
                regfile_8 <= alu_out;
              end else begin
                regfile_8 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h8 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_8 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_8 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_8 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_8 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_8 <= _T_336;
                            end else begin
                              regfile_8 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_8 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h8 == _T_150) begin
                  if (_T_304) begin
                    regfile_8 <= pc_a4;
                  end else begin
                    regfile_8 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h8 == _T_150) begin
                    if (_T_304) begin
                      regfile_8 <= csr_rdata;
                    end else begin
                      regfile_8 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h8 == _T_150) begin
            if (_T_304) begin
              regfile_8 <= alu_out;
            end else begin
              regfile_8 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h8 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_8 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_8 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_8 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_8 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_8 <= _T_336;
                          end else begin
                            regfile_8 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_8 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h8 == _T_150) begin
                if (_T_304) begin
                  regfile_8 <= pc_a4;
                end else begin
                  regfile_8 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h8 == _T_150) begin
                  if (_T_304) begin
                    regfile_8 <= csr_rdata;
                  end else begin
                    regfile_8 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h9 == io_ddpath_addr) begin
        regfile_9 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h9 == _T_150) begin
              if (_T_304) begin
                regfile_9 <= alu_out;
              end else begin
                regfile_9 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h9 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_9 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_9 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_9 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_9 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_9 <= _T_336;
                            end else begin
                              regfile_9 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_9 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h9 == _T_150) begin
                  if (_T_304) begin
                    regfile_9 <= pc_a4;
                  end else begin
                    regfile_9 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h9 == _T_150) begin
                    if (_T_304) begin
                      regfile_9 <= csr_rdata;
                    end else begin
                      regfile_9 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h9 == _T_150) begin
            if (_T_304) begin
              regfile_9 <= alu_out;
            end else begin
              regfile_9 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h9 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_9 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_9 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_9 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_9 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_9 <= _T_336;
                          end else begin
                            regfile_9 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_9 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h9 == _T_150) begin
                if (_T_304) begin
                  regfile_9 <= pc_a4;
                end else begin
                  regfile_9 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h9 == _T_150) begin
                  if (_T_304) begin
                    regfile_9 <= csr_rdata;
                  end else begin
                    regfile_9 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'ha == io_ddpath_addr) begin
        regfile_10 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'ha == _T_150) begin
              if (_T_304) begin
                regfile_10 <= alu_out;
              end else begin
                regfile_10 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'ha == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_10 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_10 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_10 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_10 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_10 <= _T_336;
                            end else begin
                              regfile_10 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_10 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'ha == _T_150) begin
                  if (_T_304) begin
                    regfile_10 <= pc_a4;
                  end else begin
                    regfile_10 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'ha == _T_150) begin
                    if (_T_304) begin
                      regfile_10 <= csr_rdata;
                    end else begin
                      regfile_10 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'ha == _T_150) begin
            if (_T_304) begin
              regfile_10 <= alu_out;
            end else begin
              regfile_10 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'ha == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_10 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_10 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_10 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_10 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_10 <= _T_336;
                          end else begin
                            regfile_10 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_10 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'ha == _T_150) begin
                if (_T_304) begin
                  regfile_10 <= pc_a4;
                end else begin
                  regfile_10 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'ha == _T_150) begin
                  if (_T_304) begin
                    regfile_10 <= csr_rdata;
                  end else begin
                    regfile_10 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'hb == io_ddpath_addr) begin
        regfile_11 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'hb == _T_150) begin
              if (_T_304) begin
                regfile_11 <= alu_out;
              end else begin
                regfile_11 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'hb == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_11 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_11 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_11 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_11 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_11 <= _T_336;
                            end else begin
                              regfile_11 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_11 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'hb == _T_150) begin
                  if (_T_304) begin
                    regfile_11 <= pc_a4;
                  end else begin
                    regfile_11 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'hb == _T_150) begin
                    if (_T_304) begin
                      regfile_11 <= csr_rdata;
                    end else begin
                      regfile_11 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'hb == _T_150) begin
            if (_T_304) begin
              regfile_11 <= alu_out;
            end else begin
              regfile_11 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'hb == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_11 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_11 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_11 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_11 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_11 <= _T_336;
                          end else begin
                            regfile_11 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_11 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'hb == _T_150) begin
                if (_T_304) begin
                  regfile_11 <= pc_a4;
                end else begin
                  regfile_11 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'hb == _T_150) begin
                  if (_T_304) begin
                    regfile_11 <= csr_rdata;
                  end else begin
                    regfile_11 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'hc == io_ddpath_addr) begin
        regfile_12 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'hc == _T_150) begin
              if (_T_304) begin
                regfile_12 <= alu_out;
              end else begin
                regfile_12 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'hc == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_12 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_12 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_12 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_12 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_12 <= _T_336;
                            end else begin
                              regfile_12 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_12 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'hc == _T_150) begin
                  if (_T_304) begin
                    regfile_12 <= pc_a4;
                  end else begin
                    regfile_12 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'hc == _T_150) begin
                    if (_T_304) begin
                      regfile_12 <= csr_rdata;
                    end else begin
                      regfile_12 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'hc == _T_150) begin
            if (_T_304) begin
              regfile_12 <= alu_out;
            end else begin
              regfile_12 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'hc == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_12 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_12 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_12 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_12 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_12 <= _T_336;
                          end else begin
                            regfile_12 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_12 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'hc == _T_150) begin
                if (_T_304) begin
                  regfile_12 <= pc_a4;
                end else begin
                  regfile_12 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'hc == _T_150) begin
                  if (_T_304) begin
                    regfile_12 <= csr_rdata;
                  end else begin
                    regfile_12 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'hd == io_ddpath_addr) begin
        regfile_13 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'hd == _T_150) begin
              if (_T_304) begin
                regfile_13 <= alu_out;
              end else begin
                regfile_13 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'hd == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_13 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_13 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_13 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_13 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_13 <= _T_336;
                            end else begin
                              regfile_13 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_13 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'hd == _T_150) begin
                  if (_T_304) begin
                    regfile_13 <= pc_a4;
                  end else begin
                    regfile_13 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'hd == _T_150) begin
                    if (_T_304) begin
                      regfile_13 <= csr_rdata;
                    end else begin
                      regfile_13 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'hd == _T_150) begin
            if (_T_304) begin
              regfile_13 <= alu_out;
            end else begin
              regfile_13 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'hd == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_13 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_13 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_13 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_13 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_13 <= _T_336;
                          end else begin
                            regfile_13 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_13 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'hd == _T_150) begin
                if (_T_304) begin
                  regfile_13 <= pc_a4;
                end else begin
                  regfile_13 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'hd == _T_150) begin
                  if (_T_304) begin
                    regfile_13 <= csr_rdata;
                  end else begin
                    regfile_13 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'he == io_ddpath_addr) begin
        regfile_14 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'he == _T_150) begin
              if (_T_304) begin
                regfile_14 <= alu_out;
              end else begin
                regfile_14 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'he == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_14 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_14 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_14 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_14 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_14 <= _T_336;
                            end else begin
                              regfile_14 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_14 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'he == _T_150) begin
                  if (_T_304) begin
                    regfile_14 <= pc_a4;
                  end else begin
                    regfile_14 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'he == _T_150) begin
                    if (_T_304) begin
                      regfile_14 <= csr_rdata;
                    end else begin
                      regfile_14 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'he == _T_150) begin
            if (_T_304) begin
              regfile_14 <= alu_out;
            end else begin
              regfile_14 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'he == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_14 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_14 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_14 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_14 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_14 <= _T_336;
                          end else begin
                            regfile_14 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_14 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'he == _T_150) begin
                if (_T_304) begin
                  regfile_14 <= pc_a4;
                end else begin
                  regfile_14 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'he == _T_150) begin
                  if (_T_304) begin
                    regfile_14 <= csr_rdata;
                  end else begin
                    regfile_14 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'hf == io_ddpath_addr) begin
        regfile_15 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'hf == _T_150) begin
              if (_T_304) begin
                regfile_15 <= alu_out;
              end else begin
                regfile_15 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'hf == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_15 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_15 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_15 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_15 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_15 <= _T_336;
                            end else begin
                              regfile_15 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_15 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'hf == _T_150) begin
                  if (_T_304) begin
                    regfile_15 <= pc_a4;
                  end else begin
                    regfile_15 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'hf == _T_150) begin
                    if (_T_304) begin
                      regfile_15 <= csr_rdata;
                    end else begin
                      regfile_15 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'hf == _T_150) begin
            if (_T_304) begin
              regfile_15 <= alu_out;
            end else begin
              regfile_15 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'hf == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_15 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_15 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_15 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_15 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_15 <= _T_336;
                          end else begin
                            regfile_15 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_15 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'hf == _T_150) begin
                if (_T_304) begin
                  regfile_15 <= pc_a4;
                end else begin
                  regfile_15 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'hf == _T_150) begin
                  if (_T_304) begin
                    regfile_15 <= csr_rdata;
                  end else begin
                    regfile_15 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h10 == io_ddpath_addr) begin
        regfile_16 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h10 == _T_150) begin
              if (_T_304) begin
                regfile_16 <= alu_out;
              end else begin
                regfile_16 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h10 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_16 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_16 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_16 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_16 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_16 <= _T_336;
                            end else begin
                              regfile_16 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_16 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h10 == _T_150) begin
                  if (_T_304) begin
                    regfile_16 <= pc_a4;
                  end else begin
                    regfile_16 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h10 == _T_150) begin
                    if (_T_304) begin
                      regfile_16 <= csr_rdata;
                    end else begin
                      regfile_16 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h10 == _T_150) begin
            if (_T_304) begin
              regfile_16 <= alu_out;
            end else begin
              regfile_16 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h10 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_16 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_16 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_16 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_16 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_16 <= _T_336;
                          end else begin
                            regfile_16 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_16 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h10 == _T_150) begin
                if (_T_304) begin
                  regfile_16 <= pc_a4;
                end else begin
                  regfile_16 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h10 == _T_150) begin
                  if (_T_304) begin
                    regfile_16 <= csr_rdata;
                  end else begin
                    regfile_16 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h11 == io_ddpath_addr) begin
        regfile_17 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h11 == _T_150) begin
              if (_T_304) begin
                regfile_17 <= alu_out;
              end else begin
                regfile_17 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h11 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_17 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_17 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_17 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_17 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_17 <= _T_336;
                            end else begin
                              regfile_17 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_17 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h11 == _T_150) begin
                  if (_T_304) begin
                    regfile_17 <= pc_a4;
                  end else begin
                    regfile_17 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h11 == _T_150) begin
                    if (_T_304) begin
                      regfile_17 <= csr_rdata;
                    end else begin
                      regfile_17 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h11 == _T_150) begin
            if (_T_304) begin
              regfile_17 <= alu_out;
            end else begin
              regfile_17 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h11 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_17 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_17 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_17 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_17 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_17 <= _T_336;
                          end else begin
                            regfile_17 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_17 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h11 == _T_150) begin
                if (_T_304) begin
                  regfile_17 <= pc_a4;
                end else begin
                  regfile_17 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h11 == _T_150) begin
                  if (_T_304) begin
                    regfile_17 <= csr_rdata;
                  end else begin
                    regfile_17 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h12 == io_ddpath_addr) begin
        regfile_18 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h12 == _T_150) begin
              if (_T_304) begin
                regfile_18 <= alu_out;
              end else begin
                regfile_18 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h12 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_18 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_18 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_18 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_18 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_18 <= _T_336;
                            end else begin
                              regfile_18 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_18 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h12 == _T_150) begin
                  if (_T_304) begin
                    regfile_18 <= pc_a4;
                  end else begin
                    regfile_18 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h12 == _T_150) begin
                    if (_T_304) begin
                      regfile_18 <= csr_rdata;
                    end else begin
                      regfile_18 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h12 == _T_150) begin
            if (_T_304) begin
              regfile_18 <= alu_out;
            end else begin
              regfile_18 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h12 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_18 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_18 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_18 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_18 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_18 <= _T_336;
                          end else begin
                            regfile_18 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_18 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h12 == _T_150) begin
                if (_T_304) begin
                  regfile_18 <= pc_a4;
                end else begin
                  regfile_18 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h12 == _T_150) begin
                  if (_T_304) begin
                    regfile_18 <= csr_rdata;
                  end else begin
                    regfile_18 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h13 == io_ddpath_addr) begin
        regfile_19 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h13 == _T_150) begin
              if (_T_304) begin
                regfile_19 <= alu_out;
              end else begin
                regfile_19 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h13 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_19 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_19 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_19 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_19 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_19 <= _T_336;
                            end else begin
                              regfile_19 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_19 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h13 == _T_150) begin
                  if (_T_304) begin
                    regfile_19 <= pc_a4;
                  end else begin
                    regfile_19 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h13 == _T_150) begin
                    if (_T_304) begin
                      regfile_19 <= csr_rdata;
                    end else begin
                      regfile_19 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h13 == _T_150) begin
            if (_T_304) begin
              regfile_19 <= alu_out;
            end else begin
              regfile_19 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h13 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_19 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_19 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_19 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_19 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_19 <= _T_336;
                          end else begin
                            regfile_19 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_19 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h13 == _T_150) begin
                if (_T_304) begin
                  regfile_19 <= pc_a4;
                end else begin
                  regfile_19 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h13 == _T_150) begin
                  if (_T_304) begin
                    regfile_19 <= csr_rdata;
                  end else begin
                    regfile_19 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h14 == io_ddpath_addr) begin
        regfile_20 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h14 == _T_150) begin
              if (_T_304) begin
                regfile_20 <= alu_out;
              end else begin
                regfile_20 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h14 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_20 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_20 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_20 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_20 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_20 <= _T_336;
                            end else begin
                              regfile_20 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_20 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h14 == _T_150) begin
                  if (_T_304) begin
                    regfile_20 <= pc_a4;
                  end else begin
                    regfile_20 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h14 == _T_150) begin
                    if (_T_304) begin
                      regfile_20 <= csr_rdata;
                    end else begin
                      regfile_20 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h14 == _T_150) begin
            if (_T_304) begin
              regfile_20 <= alu_out;
            end else begin
              regfile_20 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h14 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_20 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_20 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_20 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_20 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_20 <= _T_336;
                          end else begin
                            regfile_20 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_20 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h14 == _T_150) begin
                if (_T_304) begin
                  regfile_20 <= pc_a4;
                end else begin
                  regfile_20 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h14 == _T_150) begin
                  if (_T_304) begin
                    regfile_20 <= csr_rdata;
                  end else begin
                    regfile_20 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h15 == io_ddpath_addr) begin
        regfile_21 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h15 == _T_150) begin
              if (_T_304) begin
                regfile_21 <= alu_out;
              end else begin
                regfile_21 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h15 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_21 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_21 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_21 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_21 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_21 <= _T_336;
                            end else begin
                              regfile_21 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_21 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h15 == _T_150) begin
                  if (_T_304) begin
                    regfile_21 <= pc_a4;
                  end else begin
                    regfile_21 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h15 == _T_150) begin
                    if (_T_304) begin
                      regfile_21 <= csr_rdata;
                    end else begin
                      regfile_21 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h15 == _T_150) begin
            if (_T_304) begin
              regfile_21 <= alu_out;
            end else begin
              regfile_21 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h15 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_21 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_21 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_21 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_21 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_21 <= _T_336;
                          end else begin
                            regfile_21 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_21 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h15 == _T_150) begin
                if (_T_304) begin
                  regfile_21 <= pc_a4;
                end else begin
                  regfile_21 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h15 == _T_150) begin
                  if (_T_304) begin
                    regfile_21 <= csr_rdata;
                  end else begin
                    regfile_21 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h16 == io_ddpath_addr) begin
        regfile_22 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h16 == _T_150) begin
              if (_T_304) begin
                regfile_22 <= alu_out;
              end else begin
                regfile_22 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h16 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_22 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_22 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_22 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_22 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_22 <= _T_336;
                            end else begin
                              regfile_22 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_22 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h16 == _T_150) begin
                  if (_T_304) begin
                    regfile_22 <= pc_a4;
                  end else begin
                    regfile_22 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h16 == _T_150) begin
                    if (_T_304) begin
                      regfile_22 <= csr_rdata;
                    end else begin
                      regfile_22 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h16 == _T_150) begin
            if (_T_304) begin
              regfile_22 <= alu_out;
            end else begin
              regfile_22 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h16 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_22 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_22 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_22 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_22 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_22 <= _T_336;
                          end else begin
                            regfile_22 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_22 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h16 == _T_150) begin
                if (_T_304) begin
                  regfile_22 <= pc_a4;
                end else begin
                  regfile_22 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h16 == _T_150) begin
                  if (_T_304) begin
                    regfile_22 <= csr_rdata;
                  end else begin
                    regfile_22 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h17 == io_ddpath_addr) begin
        regfile_23 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h17 == _T_150) begin
              if (_T_304) begin
                regfile_23 <= alu_out;
              end else begin
                regfile_23 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h17 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_23 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_23 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_23 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_23 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_23 <= _T_336;
                            end else begin
                              regfile_23 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_23 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h17 == _T_150) begin
                  if (_T_304) begin
                    regfile_23 <= pc_a4;
                  end else begin
                    regfile_23 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h17 == _T_150) begin
                    if (_T_304) begin
                      regfile_23 <= csr_rdata;
                    end else begin
                      regfile_23 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h17 == _T_150) begin
            if (_T_304) begin
              regfile_23 <= alu_out;
            end else begin
              regfile_23 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h17 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_23 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_23 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_23 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_23 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_23 <= _T_336;
                          end else begin
                            regfile_23 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_23 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h17 == _T_150) begin
                if (_T_304) begin
                  regfile_23 <= pc_a4;
                end else begin
                  regfile_23 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h17 == _T_150) begin
                  if (_T_304) begin
                    regfile_23 <= csr_rdata;
                  end else begin
                    regfile_23 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h18 == io_ddpath_addr) begin
        regfile_24 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h18 == _T_150) begin
              if (_T_304) begin
                regfile_24 <= alu_out;
              end else begin
                regfile_24 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h18 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_24 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_24 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_24 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_24 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_24 <= _T_336;
                            end else begin
                              regfile_24 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_24 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h18 == _T_150) begin
                  if (_T_304) begin
                    regfile_24 <= pc_a4;
                  end else begin
                    regfile_24 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h18 == _T_150) begin
                    if (_T_304) begin
                      regfile_24 <= csr_rdata;
                    end else begin
                      regfile_24 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h18 == _T_150) begin
            if (_T_304) begin
              regfile_24 <= alu_out;
            end else begin
              regfile_24 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h18 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_24 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_24 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_24 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_24 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_24 <= _T_336;
                          end else begin
                            regfile_24 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_24 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h18 == _T_150) begin
                if (_T_304) begin
                  regfile_24 <= pc_a4;
                end else begin
                  regfile_24 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h18 == _T_150) begin
                  if (_T_304) begin
                    regfile_24 <= csr_rdata;
                  end else begin
                    regfile_24 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h19 == io_ddpath_addr) begin
        regfile_25 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h19 == _T_150) begin
              if (_T_304) begin
                regfile_25 <= alu_out;
              end else begin
                regfile_25 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h19 == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_25 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_25 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_25 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_25 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_25 <= _T_336;
                            end else begin
                              regfile_25 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_25 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h19 == _T_150) begin
                  if (_T_304) begin
                    regfile_25 <= pc_a4;
                  end else begin
                    regfile_25 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h19 == _T_150) begin
                    if (_T_304) begin
                      regfile_25 <= csr_rdata;
                    end else begin
                      regfile_25 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h19 == _T_150) begin
            if (_T_304) begin
              regfile_25 <= alu_out;
            end else begin
              regfile_25 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h19 == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_25 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_25 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_25 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_25 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_25 <= _T_336;
                          end else begin
                            regfile_25 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_25 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h19 == _T_150) begin
                if (_T_304) begin
                  regfile_25 <= pc_a4;
                end else begin
                  regfile_25 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h19 == _T_150) begin
                  if (_T_304) begin
                    regfile_25 <= csr_rdata;
                  end else begin
                    regfile_25 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h1a == io_ddpath_addr) begin
        regfile_26 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h1a == _T_150) begin
              if (_T_304) begin
                regfile_26 <= alu_out;
              end else begin
                regfile_26 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h1a == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_26 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_26 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_26 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_26 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_26 <= _T_336;
                            end else begin
                              regfile_26 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_26 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h1a == _T_150) begin
                  if (_T_304) begin
                    regfile_26 <= pc_a4;
                  end else begin
                    regfile_26 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h1a == _T_150) begin
                    if (_T_304) begin
                      regfile_26 <= csr_rdata;
                    end else begin
                      regfile_26 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h1a == _T_150) begin
            if (_T_304) begin
              regfile_26 <= alu_out;
            end else begin
              regfile_26 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h1a == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_26 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_26 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_26 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_26 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_26 <= _T_336;
                          end else begin
                            regfile_26 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_26 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h1a == _T_150) begin
                if (_T_304) begin
                  regfile_26 <= pc_a4;
                end else begin
                  regfile_26 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h1a == _T_150) begin
                  if (_T_304) begin
                    regfile_26 <= csr_rdata;
                  end else begin
                    regfile_26 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h1b == io_ddpath_addr) begin
        regfile_27 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h1b == _T_150) begin
              if (_T_304) begin
                regfile_27 <= alu_out;
              end else begin
                regfile_27 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h1b == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_27 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_27 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_27 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_27 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_27 <= _T_336;
                            end else begin
                              regfile_27 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_27 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h1b == _T_150) begin
                  if (_T_304) begin
                    regfile_27 <= pc_a4;
                  end else begin
                    regfile_27 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h1b == _T_150) begin
                    if (_T_304) begin
                      regfile_27 <= csr_rdata;
                    end else begin
                      regfile_27 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h1b == _T_150) begin
            if (_T_304) begin
              regfile_27 <= alu_out;
            end else begin
              regfile_27 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h1b == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_27 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_27 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_27 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_27 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_27 <= _T_336;
                          end else begin
                            regfile_27 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_27 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h1b == _T_150) begin
                if (_T_304) begin
                  regfile_27 <= pc_a4;
                end else begin
                  regfile_27 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h1b == _T_150) begin
                  if (_T_304) begin
                    regfile_27 <= csr_rdata;
                  end else begin
                    regfile_27 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h1c == io_ddpath_addr) begin
        regfile_28 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h1c == _T_150) begin
              if (_T_304) begin
                regfile_28 <= alu_out;
              end else begin
                regfile_28 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h1c == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_28 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_28 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_28 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_28 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_28 <= _T_336;
                            end else begin
                              regfile_28 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_28 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h1c == _T_150) begin
                  if (_T_304) begin
                    regfile_28 <= pc_a4;
                  end else begin
                    regfile_28 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h1c == _T_150) begin
                    if (_T_304) begin
                      regfile_28 <= csr_rdata;
                    end else begin
                      regfile_28 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h1c == _T_150) begin
            if (_T_304) begin
              regfile_28 <= alu_out;
            end else begin
              regfile_28 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h1c == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_28 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_28 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_28 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_28 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_28 <= _T_336;
                          end else begin
                            regfile_28 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_28 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h1c == _T_150) begin
                if (_T_304) begin
                  regfile_28 <= pc_a4;
                end else begin
                  regfile_28 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h1c == _T_150) begin
                  if (_T_304) begin
                    regfile_28 <= csr_rdata;
                  end else begin
                    regfile_28 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h1d == io_ddpath_addr) begin
        regfile_29 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h1d == _T_150) begin
              if (_T_304) begin
                regfile_29 <= alu_out;
              end else begin
                regfile_29 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h1d == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_29 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_29 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_29 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_29 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_29 <= _T_336;
                            end else begin
                              regfile_29 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_29 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h1d == _T_150) begin
                  if (_T_304) begin
                    regfile_29 <= pc_a4;
                  end else begin
                    regfile_29 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h1d == _T_150) begin
                    if (_T_304) begin
                      regfile_29 <= csr_rdata;
                    end else begin
                      regfile_29 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h1d == _T_150) begin
            if (_T_304) begin
              regfile_29 <= alu_out;
            end else begin
              regfile_29 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h1d == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_29 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_29 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_29 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_29 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_29 <= _T_336;
                          end else begin
                            regfile_29 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_29 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h1d == _T_150) begin
                if (_T_304) begin
                  regfile_29 <= pc_a4;
                end else begin
                  regfile_29 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h1d == _T_150) begin
                  if (_T_304) begin
                    regfile_29 <= csr_rdata;
                  end else begin
                    regfile_29 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h1e == io_ddpath_addr) begin
        regfile_30 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h1e == _T_150) begin
              if (_T_304) begin
                regfile_30 <= alu_out;
              end else begin
                regfile_30 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h1e == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_30 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_30 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_30 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_30 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_30 <= _T_336;
                            end else begin
                              regfile_30 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_30 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h1e == _T_150) begin
                  if (_T_304) begin
                    regfile_30 <= pc_a4;
                  end else begin
                    regfile_30 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h1e == _T_150) begin
                    if (_T_304) begin
                      regfile_30 <= csr_rdata;
                    end else begin
                      regfile_30 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h1e == _T_150) begin
            if (_T_304) begin
              regfile_30 <= alu_out;
            end else begin
              regfile_30 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h1e == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_30 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_30 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_30 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_30 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_30 <= _T_336;
                          end else begin
                            regfile_30 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_30 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h1e == _T_150) begin
                if (_T_304) begin
                  regfile_30 <= pc_a4;
                end else begin
                  regfile_30 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h1e == _T_150) begin
                  if (_T_304) begin
                    regfile_30 <= csr_rdata;
                  end else begin
                    regfile_30 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_ddpath_valid) begin
      if (5'h1f == io_ddpath_addr) begin
        regfile_31 <= io_ddpath_wdata;
      end else begin
        if (io_c2d_reg_wren) begin
          if (_T_301) begin
            if (5'h1f == _T_150) begin
              if (_T_304) begin
                regfile_31 <= alu_out;
              end else begin
                regfile_31 <= 32'h0;
              end
            end
          end else begin
            if (_T_307) begin
              if (io_dmem_resp_valid) begin
                if (5'h1f == _T_150) begin
                  if (_T_304) begin
                    if (_T_299) begin
                      regfile_31 <= _T_315;
                    end else begin
                      if (_T_297) begin
                        regfile_31 <= _T_322;
                      end else begin
                        if (_T_295) begin
                          regfile_31 <= io_dmem_resp_data;
                        end else begin
                          if (_T_293) begin
                            regfile_31 <= _T_329;
                          end else begin
                            if (_T_291) begin
                              regfile_31 <= _T_336;
                            end else begin
                              regfile_31 <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    regfile_31 <= 32'h0;
                  end
                end
              end
            end else begin
              if (_T_352) begin
                if (5'h1f == _T_150) begin
                  if (_T_304) begin
                    regfile_31 <= pc_a4;
                  end else begin
                    regfile_31 <= 32'h0;
                  end
                end
              end else begin
                if (_T_358) begin
                  if (5'h1f == _T_150) begin
                    if (_T_304) begin
                      regfile_31 <= csr_rdata;
                    end else begin
                      regfile_31 <= 32'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (io_c2d_reg_wren) begin
        if (_T_301) begin
          if (5'h1f == _T_150) begin
            if (_T_304) begin
              regfile_31 <= alu_out;
            end else begin
              regfile_31 <= 32'h0;
            end
          end
        end else begin
          if (_T_307) begin
            if (io_dmem_resp_valid) begin
              if (5'h1f == _T_150) begin
                if (_T_304) begin
                  if (_T_299) begin
                    regfile_31 <= _T_315;
                  end else begin
                    if (_T_297) begin
                      regfile_31 <= _T_322;
                    end else begin
                      if (_T_295) begin
                        regfile_31 <= io_dmem_resp_data;
                      end else begin
                        if (_T_293) begin
                          regfile_31 <= _T_329;
                        end else begin
                          if (_T_291) begin
                            regfile_31 <= _T_336;
                          end else begin
                            regfile_31 <= 32'h0;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  regfile_31 <= 32'h0;
                end
              end
            end
          end else begin
            if (_T_352) begin
              if (5'h1f == _T_150) begin
                if (_T_304) begin
                  regfile_31 <= pc_a4;
                end else begin
                  regfile_31 <= 32'h0;
                end
              end
            end else begin
              if (_T_358) begin
                if (5'h1f == _T_150) begin
                  if (_T_304) begin
                    regfile_31 <= csr_rdata;
                  end else begin
                    regfile_31 <= 32'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module rvcore( // @[:@3766.2]
  input         clock, // @[:@3767.4]
  input         reset, // @[:@3768.4]
  output [31:0] io_imem_req_addr, // @[:@3769.4]
  output        io_imem_req_valid, // @[:@3769.4]
  input  [31:0] io_imem_resp_data, // @[:@3769.4]
  input         io_imem_resp_valid, // @[:@3769.4]
  output [31:0] io_dmem_req_addr, // @[:@3769.4]
  output [31:0] io_dmem_req_data, // @[:@3769.4]
  output        io_dmem_req_mfunc, // @[:@3769.4]
  output [1:0]  io_dmem_req_mtype, // @[:@3769.4]
  output        io_dmem_req_valid, // @[:@3769.4]
  input         io_dmem_req_ready, // @[:@3769.4]
  input  [31:0] io_dmem_resp_data, // @[:@3769.4]
  input         io_dmem_resp_valid, // @[:@3769.4]
  input  [4:0]  io_ddpath_addr, // @[:@3769.4]
  input  [31:0] io_ddpath_wdata, // @[:@3769.4]
  input         io_ddpath_valid, // @[:@3769.4]
  output [31:0] io_ddpath_rdata // @[:@3769.4]
);
  wire [31:0] cpath_io_d2c_inst; // @[rvcore.scala 28:23:@3771.4]
  wire  cpath_io_d2c_dexcp; // @[rvcore.scala 28:23:@3771.4]
  wire [3:0] cpath_io_c2d_alu_func; // @[rvcore.scala 28:23:@3771.4]
  wire [2:0] cpath_io_c2d_op2_sel; // @[rvcore.scala 28:23:@3771.4]
  wire  cpath_io_c2d_reg_wren; // @[rvcore.scala 28:23:@3771.4]
  wire  cpath_io_c2d_mem_wren; // @[rvcore.scala 28:23:@3771.4]
  wire  cpath_io_c2d_mem_en; // @[rvcore.scala 28:23:@3771.4]
  wire [1:0] cpath_io_c2d_wb_sel; // @[rvcore.scala 28:23:@3771.4]
  wire [2:0] cpath_io_c2d_mem_type; // @[rvcore.scala 28:23:@3771.4]
  wire [1:0] cpath_io_c2d_pc_sel; // @[rvcore.scala 28:23:@3771.4]
  wire [2:0] cpath_io_c2d_br_sel; // @[rvcore.scala 28:23:@3771.4]
  wire [1:0] cpath_io_c2d_op1_sel; // @[rvcore.scala 28:23:@3771.4]
  wire [2:0] cpath_io_c2d_csr_cmd; // @[rvcore.scala 28:23:@3771.4]
  wire  cpath_io_c2d_cexcp; // @[rvcore.scala 28:23:@3771.4]
  wire [3:0] cpath_io_c2d_ccause; // @[rvcore.scala 28:23:@3771.4]
  wire  dpath_clock; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_reset; // @[rvcore.scala 29:23:@3774.4]
  wire [31:0] dpath_io_imem_req_addr; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_imem_req_valid; // @[rvcore.scala 29:23:@3774.4]
  wire [31:0] dpath_io_imem_resp_data; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_imem_resp_valid; // @[rvcore.scala 29:23:@3774.4]
  wire [31:0] dpath_io_dmem_req_addr; // @[rvcore.scala 29:23:@3774.4]
  wire [31:0] dpath_io_dmem_req_data; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_dmem_req_mfunc; // @[rvcore.scala 29:23:@3774.4]
  wire [1:0] dpath_io_dmem_req_mtype; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_dmem_req_valid; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_dmem_req_ready; // @[rvcore.scala 29:23:@3774.4]
  wire [31:0] dpath_io_dmem_resp_data; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_dmem_resp_valid; // @[rvcore.scala 29:23:@3774.4]
  wire [31:0] dpath_io_d2c_inst; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_d2c_dexcp; // @[rvcore.scala 29:23:@3774.4]
  wire [3:0] dpath_io_c2d_alu_func; // @[rvcore.scala 29:23:@3774.4]
  wire [2:0] dpath_io_c2d_op2_sel; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_c2d_reg_wren; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_c2d_mem_wren; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_c2d_mem_en; // @[rvcore.scala 29:23:@3774.4]
  wire [1:0] dpath_io_c2d_wb_sel; // @[rvcore.scala 29:23:@3774.4]
  wire [2:0] dpath_io_c2d_mem_type; // @[rvcore.scala 29:23:@3774.4]
  wire [1:0] dpath_io_c2d_pc_sel; // @[rvcore.scala 29:23:@3774.4]
  wire [2:0] dpath_io_c2d_br_sel; // @[rvcore.scala 29:23:@3774.4]
  wire [1:0] dpath_io_c2d_op1_sel; // @[rvcore.scala 29:23:@3774.4]
  wire [2:0] dpath_io_c2d_csr_cmd; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_c2d_cexcp; // @[rvcore.scala 29:23:@3774.4]
  wire [3:0] dpath_io_c2d_ccause; // @[rvcore.scala 29:23:@3774.4]
  wire [4:0] dpath_io_ddpath_addr; // @[rvcore.scala 29:23:@3774.4]
  wire [31:0] dpath_io_ddpath_wdata; // @[rvcore.scala 29:23:@3774.4]
  wire  dpath_io_ddpath_valid; // @[rvcore.scala 29:23:@3774.4]
  wire [31:0] dpath_io_ddpath_rdata; // @[rvcore.scala 29:23:@3774.4]
  rvcpath cpath ( // @[rvcore.scala 28:23:@3771.4]
    .io_d2c_inst(cpath_io_d2c_inst),
    .io_d2c_dexcp(cpath_io_d2c_dexcp),
    .io_c2d_alu_func(cpath_io_c2d_alu_func),
    .io_c2d_op2_sel(cpath_io_c2d_op2_sel),
    .io_c2d_reg_wren(cpath_io_c2d_reg_wren),
    .io_c2d_mem_wren(cpath_io_c2d_mem_wren),
    .io_c2d_mem_en(cpath_io_c2d_mem_en),
    .io_c2d_wb_sel(cpath_io_c2d_wb_sel),
    .io_c2d_mem_type(cpath_io_c2d_mem_type),
    .io_c2d_pc_sel(cpath_io_c2d_pc_sel),
    .io_c2d_br_sel(cpath_io_c2d_br_sel),
    .io_c2d_op1_sel(cpath_io_c2d_op1_sel),
    .io_c2d_csr_cmd(cpath_io_c2d_csr_cmd),
    .io_c2d_cexcp(cpath_io_c2d_cexcp),
    .io_c2d_ccause(cpath_io_c2d_ccause)
  );
  rvdpath dpath ( // @[rvcore.scala 29:23:@3774.4]
    .clock(dpath_clock),
    .reset(dpath_reset),
    .io_imem_req_addr(dpath_io_imem_req_addr),
    .io_imem_req_valid(dpath_io_imem_req_valid),
    .io_imem_resp_data(dpath_io_imem_resp_data),
    .io_imem_resp_valid(dpath_io_imem_resp_valid),
    .io_dmem_req_addr(dpath_io_dmem_req_addr),
    .io_dmem_req_data(dpath_io_dmem_req_data),
    .io_dmem_req_mfunc(dpath_io_dmem_req_mfunc),
    .io_dmem_req_mtype(dpath_io_dmem_req_mtype),
    .io_dmem_req_valid(dpath_io_dmem_req_valid),
    .io_dmem_req_ready(dpath_io_dmem_req_ready),
    .io_dmem_resp_data(dpath_io_dmem_resp_data),
    .io_dmem_resp_valid(dpath_io_dmem_resp_valid),
    .io_d2c_inst(dpath_io_d2c_inst),
    .io_d2c_dexcp(dpath_io_d2c_dexcp),
    .io_c2d_alu_func(dpath_io_c2d_alu_func),
    .io_c2d_op2_sel(dpath_io_c2d_op2_sel),
    .io_c2d_reg_wren(dpath_io_c2d_reg_wren),
    .io_c2d_mem_wren(dpath_io_c2d_mem_wren),
    .io_c2d_mem_en(dpath_io_c2d_mem_en),
    .io_c2d_wb_sel(dpath_io_c2d_wb_sel),
    .io_c2d_mem_type(dpath_io_c2d_mem_type),
    .io_c2d_pc_sel(dpath_io_c2d_pc_sel),
    .io_c2d_br_sel(dpath_io_c2d_br_sel),
    .io_c2d_op1_sel(dpath_io_c2d_op1_sel),
    .io_c2d_csr_cmd(dpath_io_c2d_csr_cmd),
    .io_c2d_cexcp(dpath_io_c2d_cexcp),
    .io_c2d_ccause(dpath_io_c2d_ccause),
    .io_ddpath_addr(dpath_io_ddpath_addr),
    .io_ddpath_wdata(dpath_io_ddpath_wdata),
    .io_ddpath_valid(dpath_io_ddpath_valid),
    .io_ddpath_rdata(dpath_io_ddpath_rdata)
  );
  assign io_imem_req_addr = dpath_io_imem_req_addr;
  assign io_imem_req_valid = dpath_io_imem_req_valid;
  assign io_dmem_req_addr = dpath_io_dmem_req_addr;
  assign io_dmem_req_data = dpath_io_dmem_req_data;
  assign io_dmem_req_mfunc = dpath_io_dmem_req_mfunc;
  assign io_dmem_req_mtype = dpath_io_dmem_req_mtype;
  assign io_dmem_req_valid = dpath_io_dmem_req_valid;
  assign io_ddpath_rdata = dpath_io_ddpath_rdata;
  assign cpath_io_d2c_inst = dpath_io_d2c_inst;
  assign cpath_io_d2c_dexcp = dpath_io_d2c_dexcp;
  assign dpath_clock = clock;
  assign dpath_reset = reset;
  assign dpath_io_imem_resp_data = io_imem_resp_data;
  assign dpath_io_imem_resp_valid = io_imem_resp_valid;
  assign dpath_io_dmem_req_ready = io_dmem_req_ready;
  assign dpath_io_dmem_resp_data = io_dmem_resp_data;
  assign dpath_io_dmem_resp_valid = io_dmem_resp_valid;
  assign dpath_io_c2d_alu_func = cpath_io_c2d_alu_func;
  assign dpath_io_c2d_op2_sel = cpath_io_c2d_op2_sel;
  assign dpath_io_c2d_reg_wren = cpath_io_c2d_reg_wren;
  assign dpath_io_c2d_mem_wren = cpath_io_c2d_mem_wren;
  assign dpath_io_c2d_mem_en = cpath_io_c2d_mem_en;
  assign dpath_io_c2d_wb_sel = cpath_io_c2d_wb_sel;
  assign dpath_io_c2d_mem_type = cpath_io_c2d_mem_type;
  assign dpath_io_c2d_pc_sel = cpath_io_c2d_pc_sel;
  assign dpath_io_c2d_br_sel = cpath_io_c2d_br_sel;
  assign dpath_io_c2d_op1_sel = cpath_io_c2d_op1_sel;
  assign dpath_io_c2d_csr_cmd = cpath_io_c2d_csr_cmd;
  assign dpath_io_c2d_cexcp = cpath_io_c2d_cexcp;
  assign dpath_io_c2d_ccause = cpath_io_c2d_ccause;
  assign dpath_io_ddpath_addr = io_ddpath_addr;
  assign dpath_io_ddpath_wdata = io_ddpath_wdata;
  assign dpath_io_ddpath_valid = io_ddpath_valid;
endmodule
module rvmemarb( // @[:@3831.2]
  input         clock, // @[:@3832.4]
  input         reset, // @[:@3833.4]
  input  [31:0] io_inst_port_req_addr, // @[:@3834.4]
  input         io_inst_port_req_valid, // @[:@3834.4]
  output [31:0] io_inst_port_resp_data, // @[:@3834.4]
  output        io_inst_port_resp_valid, // @[:@3834.4]
  input  [31:0] io_data_port_req_addr, // @[:@3834.4]
  input  [31:0] io_data_port_req_data, // @[:@3834.4]
  input         io_data_port_req_mfunc, // @[:@3834.4]
  input  [1:0]  io_data_port_req_mtype, // @[:@3834.4]
  input         io_data_port_req_valid, // @[:@3834.4]
  output        io_data_port_req_ready, // @[:@3834.4]
  output [31:0] io_data_port_resp_data, // @[:@3834.4]
  output        io_data_port_resp_valid, // @[:@3834.4]
  input  [31:0] io_dm_port_req_addr, // @[:@3834.4]
  input  [31:0] io_dm_port_req_data, // @[:@3834.4]
  input         io_dm_port_req_mfunc, // @[:@3834.4]
  input         io_dm_port_req_valid, // @[:@3834.4]
  output        io_dm_port_req_ready, // @[:@3834.4]
  output [31:0] io_dm_port_resp_data, // @[:@3834.4]
  output        io_dm_port_resp_valid, // @[:@3834.4]
  output        io_ext_mem_waen, // @[:@3834.4]
  output        io_ext_mem_wden, // @[:@3834.4]
  output [31:0] io_ext_mem_waddr, // @[:@3834.4]
  output [31:0] io_ext_mem_wdata, // @[:@3834.4]
  output [3:0]  io_ext_mem_wmask, // @[:@3834.4]
  input         io_ext_mem_wardy, // @[:@3834.4]
  input         io_ext_mem_wdrdy, // @[:@3834.4]
  input         io_ext_mem_wbvld, // @[:@3834.4]
  output        io_ext_mem_raen, // @[:@3834.4]
  output        io_ext_mem_rden, // @[:@3834.4]
  output [31:0] io_ext_mem_raddr, // @[:@3834.4]
  input  [31:0] io_ext_mem_rdata, // @[:@3834.4]
  input         io_ext_mem_rardy, // @[:@3834.4]
  input         io_ext_mem_rdrdy, // @[:@3834.4]
  output        io_ext_mem_clock, // @[:@3834.4]
  output        io_ext_mem_reset // @[:@3834.4]
);
  reg [1:0] reg_stat; // @[rvmemarb.scala 164:23:@3876.4]
  reg [31:0] _RAND_0;
  reg  reg_wabusy; // @[rvmemarb.scala 166:25:@3877.4]
  reg [31:0] _RAND_1;
  reg  reg_wdbusy; // @[rvmemarb.scala 167:25:@3878.4]
  reg [31:0] _RAND_2;
  reg  reg_rabusy; // @[rvmemarb.scala 168:25:@3879.4]
  reg [31:0] _RAND_3;
  reg  reg_rdbusy; // @[rvmemarb.scala 169:25:@3880.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_dmdata; // @[rvmemarb.scala 186:25:@3895.4]
  reg [31:0] _RAND_5;
  reg  reg_dmvld; // @[rvmemarb.scala 187:24:@3896.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_ipdata; // @[rvmemarb.scala 189:25:@3897.4]
  reg [31:0] _RAND_7;
  reg  reg_ipvld; // @[rvmemarb.scala 190:24:@3898.4]
  reg [31:0] _RAND_8;
  reg [31:0] reg_dpdata; // @[rvmemarb.scala 192:25:@3899.4]
  reg [31:0] _RAND_9;
  reg  reg_dpvld; // @[rvmemarb.scala 193:24:@3900.4]
  reg [31:0] _RAND_10;
  wire  _T_147; // @[Conditional.scala 37:30:@3921.4]
  wire  _GEN_0; // @[rvmemarb.scala 243:45:@3933.14]
  wire  _GEN_1; // @[rvmemarb.scala 243:45:@3933.14]
  wire  _GEN_7; // @[rvmemarb.scala 242:46:@3932.12]
  wire  _GEN_10; // @[rvmemarb.scala 239:42:@3929.10]
  wire  _GEN_28; // @[Conditional.scala 40:58:@3925.8]
  wire  _GEN_50; // @[rvmemarb.scala 225:40:@3923.6]
  wire  _T_252; // @[Conditional.scala 37:30:@4051.6]
  wire  _T_442; // @[Conditional.scala 37:30:@4268.8]
  wire  _T_467; // @[Conditional.scala 37:30:@4336.10]
  wire  _GEN_217; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_235; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_254; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_282; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_290; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_312; // @[Conditional.scala 40:58:@3922.4]
  wire  wden; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _T_157; // @[rvmemarb.scala 252:42:@3941.14]
  wire  _GEN_3; // @[rvmemarb.scala 252:50:@3942.14]
  wire  _GEN_4; // @[rvmemarb.scala 242:46:@3932.12]
  wire  _GEN_5; // @[rvmemarb.scala 242:46:@3932.12]
  wire  _GEN_6; // @[rvmemarb.scala 242:46:@3932.12]
  wire  _GEN_9; // @[rvmemarb.scala 239:42:@3929.10]
  wire  _GEN_27; // @[Conditional.scala 40:58:@3925.8]
  wire  _GEN_49; // @[rvmemarb.scala 225:40:@3923.6]
  wire  _GEN_216; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_234; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_253; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_281; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_289; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_311; // @[Conditional.scala 40:58:@3922.4]
  wire  waen; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _T_161; // @[rvmemarb.scala 261:38:@3950.12]
  wire  _GEN_8; // @[rvmemarb.scala 261:46:@3951.12]
  wire  _GEN_11; // @[rvmemarb.scala 239:42:@3929.10]
  wire  _GEN_12; // @[rvmemarb.scala 239:42:@3929.10]
  wire  _GEN_13; // @[rvmemarb.scala 239:42:@3929.10]
  wire [7:0] _T_164; // @[rvmemarb.scala 270:41:@3957.12]
  wire [7:0] _T_199; // @[rvmemarb.scala 293:41:@3984.14]
  wire [15:0] _T_221; // @[rvmemarb.scala 306:45:@3997.14]
  wire [7:0] _T_227; // @[rvmemarb.scala 314:41:@4008.16]
  wire [7:0] _T_228; // @[rvmemarb.scala 315:41:@4009.16]
  wire [15:0] _T_240; // @[rvmemarb.scala 319:45:@4016.16]
  wire [31:0] _T_241; // @[rvmemarb.scala 319:45:@4017.16]
  wire  _T_242; // @[Conditional.scala 37:30:@4023.10]
  wire  _GEN_34; // @[Conditional.scala 40:58:@3925.8]
  wire  _GEN_56; // @[rvmemarb.scala 225:40:@3923.6]
  wire  _GEN_79; // @[rvmemarb.scala 495:44:@4180.16]
  wire  _GEN_81; // @[rvmemarb.scala 472:42:@4158.14]
  wire  _GEN_98; // @[Conditional.scala 39:67:@4155.12]
  wire  _GEN_115; // @[Conditional.scala 40:58:@4056.10]
  wire  _GEN_131; // @[rvmemarb.scala 361:40:@4053.8]
  wire  _GEN_140; // @[rvmemarb.scala 621:44:@4296.16]
  wire  _GEN_142; // @[rvmemarb.scala 598:42:@4274.14]
  wire  _GEN_163; // @[rvmemarb.scala 588:42:@4270.10]
  wire  _T_564; // @[Conditional.scala 37:30:@4453.16]
  wire  _GEN_188; // @[rvmemarb.scala 823:44:@4479.20]
  wire  _GEN_190; // @[rvmemarb.scala 800:42:@4457.18]
  wire  _GEN_204; // @[Conditional.scala 39:67:@4454.16]
  wire  _GEN_226; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_244; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_262; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_269; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_296; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_318; // @[Conditional.scala 40:58:@3922.4]
  wire  raen; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _T_245; // @[rvmemarb.scala 333:34:@4028.12]
  wire  _GEN_20; // @[rvmemarb.scala 333:42:@4029.12]
  wire [31:0] _GEN_21; // @[Conditional.scala 39:67:@4024.10]
  wire  _GEN_24; // @[Conditional.scala 39:67:@4024.10]
  wire [31:0] _GEN_25; // @[Conditional.scala 40:58:@3925.8]
  wire  _GEN_26; // @[Conditional.scala 40:58:@3925.8]
  wire  _GEN_29; // @[Conditional.scala 40:58:@3925.8]
  wire  _GEN_30; // @[Conditional.scala 40:58:@3925.8]
  wire [31:0] _GEN_31; // @[Conditional.scala 40:58:@3925.8]
  wire [3:0] _GEN_32; // @[Conditional.scala 40:58:@3925.8]
  wire [31:0] _GEN_33; // @[Conditional.scala 40:58:@3925.8]
  wire  _GEN_36; // @[Conditional.scala 40:58:@3925.8]
  wire [31:0] _GEN_42; // @[rvmemarb.scala 341:47:@4036.8]
  wire  _GEN_45; // @[rvmemarb.scala 341:47:@4036.8]
  wire [1:0] _GEN_46; // @[rvmemarb.scala 341:47:@4036.8]
  wire [31:0] _GEN_47; // @[rvmemarb.scala 225:40:@3923.6]
  wire  _GEN_48; // @[rvmemarb.scala 225:40:@3923.6]
  wire  _GEN_51; // @[rvmemarb.scala 225:40:@3923.6]
  wire  _GEN_52; // @[rvmemarb.scala 225:40:@3923.6]
  wire [31:0] _GEN_53; // @[rvmemarb.scala 225:40:@3923.6]
  wire [3:0] _GEN_54; // @[rvmemarb.scala 225:40:@3923.6]
  wire [31:0] _GEN_55; // @[rvmemarb.scala 225:40:@3923.6]
  wire  _GEN_58; // @[rvmemarb.scala 225:40:@3923.6]
  wire [1:0] _GEN_59; // @[rvmemarb.scala 225:40:@3923.6]
  wire  _GEN_71; // @[rvmemarb.scala 476:45:@4162.18]
  wire  _GEN_72; // @[rvmemarb.scala 476:45:@4162.18]
  wire  _GEN_74; // @[rvmemarb.scala 486:45:@4171.18]
  wire  _GEN_76; // @[rvmemarb.scala 475:46:@4161.16]
  wire  _GEN_78; // @[rvmemarb.scala 475:46:@4161.16]
  wire  _GEN_82; // @[rvmemarb.scala 472:42:@4158.14]
  wire  _GEN_83; // @[rvmemarb.scala 472:42:@4158.14]
  wire  _GEN_84; // @[rvmemarb.scala 472:42:@4158.14]
  wire [7:0] _T_373; // @[rvmemarb.scala 514:88:@4193.18]
  wire [31:0] _T_374; // @[Cat.scala 30:58:@4194.18]
  wire [7:0] _T_381; // @[rvmemarb.scala 515:88:@4196.18]
  wire [31:0] _T_382; // @[Cat.scala 30:58:@4197.18]
  wire [7:0] _T_389; // @[rvmemarb.scala 516:88:@4199.18]
  wire [31:0] _T_390; // @[Cat.scala 30:58:@4200.18]
  wire [7:0] _T_397; // @[rvmemarb.scala 517:88:@4202.18]
  wire [31:0] _T_398; // @[Cat.scala 30:58:@4203.18]
  wire [23:0] _T_419; // @[Cat.scala 30:58:@4222.20]
  wire [31:0] _T_420; // @[Cat.scala 30:58:@4223.20]
  wire [23:0] _T_429; // @[Cat.scala 30:58:@4227.20]
  wire [31:0] _T_430; // @[Cat.scala 30:58:@4228.20]
  wire [31:0] _GEN_92; // @[rvmemarb.scala 505:37:@4189.14]
  wire  _T_439; // @[rvmemarb.scala 551:34:@4244.16]
  wire [1:0] _GEN_94; // @[rvmemarb.scala 552:62:@4246.18]
  wire [1:0] _GEN_95; // @[rvmemarb.scala 551:57:@4245.16]
  wire [1:0] _GEN_96; // @[rvmemarb.scala 546:40:@4243.14]
  wire  _GEN_99; // @[Conditional.scala 39:67:@4155.12]
  wire  _GEN_100; // @[Conditional.scala 39:67:@4155.12]
  wire  _GEN_101; // @[Conditional.scala 39:67:@4155.12]
  wire [31:0] _GEN_103; // @[Conditional.scala 39:67:@4155.12]
  wire  _GEN_104; // @[Conditional.scala 39:67:@4155.12]
  wire [1:0] _GEN_105; // @[Conditional.scala 39:67:@4155.12]
  wire  _GEN_107; // @[Conditional.scala 40:58:@4056.10]
  wire  _GEN_116; // @[Conditional.scala 40:58:@4056.10]
  wire  _GEN_117; // @[Conditional.scala 40:58:@4056.10]
  wire  _GEN_118; // @[Conditional.scala 40:58:@4056.10]
  wire [31:0] _GEN_119; // @[Conditional.scala 40:58:@4056.10]
  wire  _GEN_120; // @[Conditional.scala 40:58:@4056.10]
  wire [1:0] _GEN_121; // @[Conditional.scala 40:58:@4056.10]
  wire  _GEN_122; // @[rvmemarb.scala 361:40:@4053.8]
  wire  _GEN_126; // @[rvmemarb.scala 361:40:@4053.8]
  wire  _GEN_127; // @[rvmemarb.scala 361:40:@4053.8]
  wire [31:0] _GEN_130; // @[rvmemarb.scala 361:40:@4053.8]
  wire  _GEN_132; // @[rvmemarb.scala 361:40:@4053.8]
  wire  _GEN_133; // @[rvmemarb.scala 361:40:@4053.8]
  wire  _GEN_134; // @[rvmemarb.scala 361:40:@4053.8]
  wire [31:0] _GEN_135; // @[rvmemarb.scala 361:40:@4053.8]
  wire  _GEN_136; // @[rvmemarb.scala 361:40:@4053.8]
  wire [1:0] _GEN_137; // @[rvmemarb.scala 361:40:@4053.8]
  wire  _GEN_144; // @[rvmemarb.scala 598:42:@4274.14]
  wire [31:0] _GEN_145; // @[rvmemarb.scala 632:37:@4305.14]
  wire  _T_463; // @[rvmemarb.scala 650:39:@4320.20]
  wire [1:0] _GEN_146; // @[rvmemarb.scala 650:64:@4321.20]
  wire [1:0] _GEN_147; // @[rvmemarb.scala 647:61:@4316.18]
  wire [1:0] _GEN_148; // @[rvmemarb.scala 643:58:@4311.16]
  wire  _GEN_149; // @[rvmemarb.scala 643:58:@4311.16]
  wire  _GEN_150; // @[rvmemarb.scala 638:40:@4309.14]
  wire [1:0] _GEN_151; // @[rvmemarb.scala 638:40:@4309.14]
  wire  _GEN_152; // @[rvmemarb.scala 638:40:@4309.14]
  wire  _GEN_164; // @[rvmemarb.scala 588:42:@4270.10]
  wire  _GEN_165; // @[rvmemarb.scala 588:42:@4270.10]
  wire  _GEN_166; // @[rvmemarb.scala 588:42:@4270.10]
  wire  _GEN_168; // @[rvmemarb.scala 588:42:@4270.10]
  wire [31:0] _GEN_169; // @[rvmemarb.scala 588:42:@4270.10]
  wire [1:0] _GEN_170; // @[rvmemarb.scala 588:42:@4270.10]
  wire  _GEN_171; // @[rvmemarb.scala 588:42:@4270.10]
  wire  _GEN_172; // @[rvmemarb.scala 588:42:@4270.10]
  wire [1:0] _T_470; // @[rvmemarb.scala 684:48:@4342.16]
  wire  _T_484; // @[Conditional.scala 37:30:@4371.16]
  wire [7:0] _T_485; // @[rvmemarb.scala 721:41:@4373.18]
  wire  _T_507; // @[Mux.scala 46:19:@4382.18]
  wire [3:0] _T_508; // @[Mux.scala 46:16:@4383.18]
  wire  _T_509; // @[Mux.scala 46:19:@4384.18]
  wire [3:0] _T_510; // @[Mux.scala 46:16:@4385.18]
  wire  _T_511; // @[Mux.scala 46:19:@4386.18]
  wire [3:0] _T_512; // @[Mux.scala 46:16:@4387.18]
  wire  _T_513; // @[Mux.scala 46:19:@4388.18]
  wire [3:0] _T_514; // @[Mux.scala 46:16:@4389.18]
  wire [15:0] _T_515; // @[rvmemarb.scala 737:45:@4390.18]
  wire [31:0] _T_517; // @[rvmemarb.scala 737:45:@4392.18]
  wire  _T_518; // @[Conditional.scala 37:30:@4397.18]
  wire [7:0] _T_520; // @[rvmemarb.scala 744:41:@4400.20]
  wire  _T_532; // @[rvmemarb.scala 749:40:@4408.20]
  wire [3:0] _T_539; // @[Mux.scala 46:16:@4410.20]
  wire  _T_540; // @[Mux.scala 46:19:@4411.20]
  wire [3:0] _T_541; // @[Mux.scala 46:16:@4412.20]
  wire [15:0] _T_542; // @[rvmemarb.scala 757:45:@4413.20]
  wire [31:0] _T_544; // @[rvmemarb.scala 757:45:@4415.20]
  wire  _T_545; // @[Conditional.scala 37:30:@4420.20]
  wire [7:0] _T_548; // @[rvmemarb.scala 765:41:@4424.22]
  wire [7:0] _T_549; // @[rvmemarb.scala 766:41:@4425.22]
  wire [15:0] _T_561; // @[rvmemarb.scala 770:45:@4432.22]
  wire [31:0] _T_562; // @[rvmemarb.scala 770:45:@4433.22]
  wire [31:0] _GEN_178; // @[Conditional.scala 39:67:@4421.20]
  wire [3:0] _GEN_179; // @[Conditional.scala 39:67:@4421.20]
  wire [31:0] _GEN_180; // @[Conditional.scala 39:67:@4398.18]
  wire [3:0] _GEN_181; // @[Conditional.scala 39:67:@4398.18]
  wire [31:0] _GEN_182; // @[Conditional.scala 40:58:@4372.16]
  wire [3:0] _GEN_183; // @[Conditional.scala 40:58:@4372.16]
  wire [1:0] _GEN_184; // @[rvmemarb.scala 783:56:@4440.18]
  wire  _GEN_185; // @[rvmemarb.scala 780:37:@4437.16]
  wire [31:0] _GEN_186; // @[rvmemarb.scala 780:37:@4437.16]
  wire [1:0] _GEN_187; // @[rvmemarb.scala 780:37:@4437.16]
  wire [31:0] _T_616; // @[Mux.scala 46:16:@4504.22]
  wire [31:0] _T_618; // @[Mux.scala 46:16:@4506.22]
  wire [31:0] _T_620; // @[Mux.scala 46:16:@4508.22]
  wire [31:0] _T_622; // @[Mux.scala 46:16:@4510.22]
  wire [31:0] _T_648; // @[Mux.scala 46:16:@4529.24]
  wire [31:0] _T_650; // @[Mux.scala 46:16:@4531.24]
  wire [31:0] _GEN_192; // @[Conditional.scala 39:67:@4537.24]
  wire [31:0] _GEN_194; // @[Conditional.scala 39:67:@4516.22]
  wire  _GEN_195; // @[Conditional.scala 39:67:@4516.22]
  wire [31:0] _GEN_196; // @[Conditional.scala 40:58:@4490.20]
  wire  _GEN_197; // @[Conditional.scala 40:58:@4490.20]
  wire [31:0] _GEN_198; // @[rvmemarb.scala 834:37:@4488.18]
  wire  _GEN_199; // @[rvmemarb.scala 834:37:@4488.18]
  wire  _GEN_200; // @[rvmemarb.scala 876:40:@4542.18]
  wire [31:0] _GEN_201; // @[rvmemarb.scala 876:40:@4542.18]
  wire [1:0] _GEN_202; // @[rvmemarb.scala 876:40:@4542.18]
  wire [31:0] _GEN_203; // @[Conditional.scala 39:67:@4454.16]
  wire  _GEN_205; // @[Conditional.scala 39:67:@4454.16]
  wire  _GEN_206; // @[Conditional.scala 39:67:@4454.16]
  wire  _GEN_207; // @[Conditional.scala 39:67:@4454.16]
  wire  _GEN_208; // @[Conditional.scala 39:67:@4454.16]
  wire [31:0] _GEN_209; // @[Conditional.scala 39:67:@4454.16]
  wire  _GEN_210; // @[Conditional.scala 39:67:@4454.16]
  wire  _GEN_211; // @[Conditional.scala 39:67:@4454.16]
  wire [31:0] _GEN_212; // @[Conditional.scala 39:67:@4454.16]
  wire [1:0] _GEN_213; // @[Conditional.scala 39:67:@4454.16]
  wire [31:0] _GEN_214; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_215; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_218; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_219; // @[Conditional.scala 40:58:@4341.14]
  wire [31:0] _GEN_220; // @[Conditional.scala 40:58:@4341.14]
  wire [3:0] _GEN_221; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_222; // @[Conditional.scala 40:58:@4341.14]
  wire [31:0] _GEN_223; // @[Conditional.scala 40:58:@4341.14]
  wire [1:0] _GEN_224; // @[Conditional.scala 40:58:@4341.14]
  wire [31:0] _GEN_225; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_227; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_228; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_229; // @[Conditional.scala 40:58:@4341.14]
  wire [31:0] _GEN_230; // @[Conditional.scala 40:58:@4341.14]
  wire  _GEN_231; // @[Conditional.scala 40:58:@4341.14]
  wire [31:0] _GEN_232; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_233; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_236; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_237; // @[rvmemarb.scala 677:42:@4339.12]
  wire [31:0] _GEN_238; // @[rvmemarb.scala 677:42:@4339.12]
  wire [3:0] _GEN_239; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_240; // @[rvmemarb.scala 677:42:@4339.12]
  wire [31:0] _GEN_241; // @[rvmemarb.scala 677:42:@4339.12]
  wire [1:0] _GEN_242; // @[rvmemarb.scala 677:42:@4339.12]
  wire [31:0] _GEN_243; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_245; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_246; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_247; // @[rvmemarb.scala 677:42:@4339.12]
  wire [31:0] _GEN_248; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_249; // @[rvmemarb.scala 677:42:@4339.12]
  wire  _GEN_250; // @[Conditional.scala 39:67:@4337.10]
  wire [31:0] _GEN_251; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_252; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_255; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_256; // @[Conditional.scala 39:67:@4337.10]
  wire [31:0] _GEN_257; // @[Conditional.scala 39:67:@4337.10]
  wire [3:0] _GEN_258; // @[Conditional.scala 39:67:@4337.10]
  wire [31:0] _GEN_259; // @[Conditional.scala 39:67:@4337.10]
  wire [1:0] _GEN_260; // @[Conditional.scala 39:67:@4337.10]
  wire [31:0] _GEN_261; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_263; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_264; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_265; // @[Conditional.scala 39:67:@4337.10]
  wire [31:0] _GEN_266; // @[Conditional.scala 39:67:@4337.10]
  wire  _GEN_267; // @[Conditional.scala 39:67:@4337.10]
  wire [31:0] _GEN_268; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_270; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_271; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_272; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_274; // @[Conditional.scala 39:67:@4269.8]
  wire [31:0] _GEN_275; // @[Conditional.scala 39:67:@4269.8]
  wire [1:0] _GEN_276; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_277; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_278; // @[Conditional.scala 39:67:@4269.8]
  wire [31:0] _GEN_279; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_280; // @[Conditional.scala 39:67:@4269.8]
  wire [31:0] _GEN_283; // @[Conditional.scala 39:67:@4269.8]
  wire [3:0] _GEN_284; // @[Conditional.scala 39:67:@4269.8]
  wire [31:0] _GEN_285; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_286; // @[Conditional.scala 39:67:@4269.8]
  wire  _GEN_287; // @[Conditional.scala 39:67:@4052.6]
  wire [31:0] _GEN_288; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_291; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_292; // @[Conditional.scala 39:67:@4052.6]
  wire [31:0] _GEN_293; // @[Conditional.scala 39:67:@4052.6]
  wire [3:0] _GEN_294; // @[Conditional.scala 39:67:@4052.6]
  wire [31:0] _GEN_295; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_297; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_298; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_299; // @[Conditional.scala 39:67:@4052.6]
  wire [31:0] _GEN_300; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_301; // @[Conditional.scala 39:67:@4052.6]
  wire [1:0] _GEN_302; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_304; // @[Conditional.scala 39:67:@4052.6]
  wire [31:0] _GEN_305; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_306; // @[Conditional.scala 39:67:@4052.6]
  wire [31:0] _GEN_307; // @[Conditional.scala 39:67:@4052.6]
  wire  _GEN_308; // @[Conditional.scala 39:67:@4052.6]
  wire [31:0] waddr; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_310; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_313; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_314; // @[Conditional.scala 40:58:@3922.4]
  wire [31:0] wdata; // @[Conditional.scala 40:58:@3922.4]
  wire [3:0] wmask; // @[Conditional.scala 40:58:@3922.4]
  wire [31:0] raddr; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_319; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_320; // @[Conditional.scala 40:58:@3922.4]
  wire [1:0] _GEN_321; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_322; // @[Conditional.scala 40:58:@3922.4]
  wire [31:0] _GEN_323; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_324; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_326; // @[Conditional.scala 40:58:@3922.4]
  wire [31:0] _GEN_327; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_328; // @[Conditional.scala 40:58:@3922.4]
  wire [31:0] _GEN_329; // @[Conditional.scala 40:58:@3922.4]
  wire  _GEN_330; // @[Conditional.scala 40:58:@3922.4]
  wire [1:0] _GEN_331; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_332; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_333; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_334; // @[rvmemarb.scala 953:26:@4584.4]
  wire  rden; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_340; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_341; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_342; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_343; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_344; // @[rvmemarb.scala 953:26:@4584.4]
  wire [31:0] _GEN_345; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_346; // @[rvmemarb.scala 953:26:@4584.4]
  wire [31:0] _GEN_347; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_348; // @[rvmemarb.scala 953:26:@4584.4]
  wire [31:0] _GEN_349; // @[rvmemarb.scala 953:26:@4584.4]
  wire  _GEN_350; // @[rvmemarb.scala 953:26:@4584.4]
  assign _T_147 = 2'h0 == reg_stat; // @[Conditional.scala 37:30:@3921.4]
  assign _GEN_0 = io_ext_mem_wbvld ? 1'h0 : reg_wabusy; // @[rvmemarb.scala 243:45:@3933.14]
  assign _GEN_1 = io_ext_mem_wbvld ? 1'h0 : reg_wdbusy; // @[rvmemarb.scala 243:45:@3933.14]
  assign _GEN_7 = reg_wdbusy ? 1'h0 : 1'h1; // @[rvmemarb.scala 242:46:@3932.12]
  assign _GEN_10 = reg_wabusy ? _GEN_7 : 1'h0; // @[rvmemarb.scala 239:42:@3929.10]
  assign _GEN_28 = io_dm_port_req_mfunc ? _GEN_10 : 1'h0; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_50 = io_dm_port_req_valid ? _GEN_28 : 1'h0; // @[rvmemarb.scala 225:40:@3923.6]
  assign _T_252 = 2'h1 == reg_stat; // @[Conditional.scala 37:30:@4051.6]
  assign _T_442 = 2'h2 == reg_stat; // @[Conditional.scala 37:30:@4268.8]
  assign _T_467 = 2'h3 == reg_stat; // @[Conditional.scala 37:30:@4336.10]
  assign _GEN_217 = io_data_port_req_mfunc ? _GEN_10 : 1'h0; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_235 = io_data_port_req_valid ? _GEN_217 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_254 = _T_467 ? _GEN_235 : 1'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_282 = _T_442 ? 1'h0 : _GEN_254; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_290 = _T_252 ? _GEN_50 : _GEN_282; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_312 = _T_147 ? _GEN_50 : _GEN_290; // @[Conditional.scala 40:58:@3922.4]
  assign wden = reset ? 1'h0 : _GEN_312; // @[rvmemarb.scala 953:26:@4584.4]
  assign _T_157 = wden & io_ext_mem_wdrdy; // @[rvmemarb.scala 252:42:@3941.14]
  assign _GEN_3 = _T_157 ? 1'h1 : reg_wdbusy; // @[rvmemarb.scala 252:50:@3942.14]
  assign _GEN_4 = reg_wdbusy ? _GEN_0 : reg_wabusy; // @[rvmemarb.scala 242:46:@3932.12]
  assign _GEN_5 = reg_wdbusy ? _GEN_1 : _GEN_3; // @[rvmemarb.scala 242:46:@3932.12]
  assign _GEN_6 = reg_wdbusy ? io_ext_mem_wbvld : 1'h0; // @[rvmemarb.scala 242:46:@3932.12]
  assign _GEN_9 = reg_wabusy ? 1'h0 : 1'h1; // @[rvmemarb.scala 239:42:@3929.10]
  assign _GEN_27 = io_dm_port_req_mfunc ? _GEN_9 : 1'h0; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_49 = io_dm_port_req_valid ? _GEN_27 : 1'h0; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_216 = io_data_port_req_mfunc ? _GEN_9 : 1'h0; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_234 = io_data_port_req_valid ? _GEN_216 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_253 = _T_467 ? _GEN_234 : 1'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_281 = _T_442 ? 1'h0 : _GEN_253; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_289 = _T_252 ? _GEN_49 : _GEN_281; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_311 = _T_147 ? _GEN_49 : _GEN_289; // @[Conditional.scala 40:58:@3922.4]
  assign waen = reset ? 1'h0 : _GEN_311; // @[rvmemarb.scala 953:26:@4584.4]
  assign _T_161 = waen & io_ext_mem_wardy; // @[rvmemarb.scala 261:38:@3950.12]
  assign _GEN_8 = _T_161 ? 1'h1 : reg_wabusy; // @[rvmemarb.scala 261:46:@3951.12]
  assign _GEN_11 = reg_wabusy ? _GEN_4 : _GEN_8; // @[rvmemarb.scala 239:42:@3929.10]
  assign _GEN_12 = reg_wabusy ? _GEN_5 : reg_wdbusy; // @[rvmemarb.scala 239:42:@3929.10]
  assign _GEN_13 = reg_wabusy ? _GEN_6 : 1'h0; // @[rvmemarb.scala 239:42:@3929.10]
  assign _T_164 = io_dm_port_req_data[7:0]; // @[rvmemarb.scala 270:41:@3957.12]
  assign _T_199 = io_dm_port_req_data[15:8]; // @[rvmemarb.scala 293:41:@3984.14]
  assign _T_221 = {_T_199,_T_164}; // @[rvmemarb.scala 306:45:@3997.14]
  assign _T_227 = io_dm_port_req_data[23:16]; // @[rvmemarb.scala 314:41:@4008.16]
  assign _T_228 = io_dm_port_req_data[31:24]; // @[rvmemarb.scala 315:41:@4009.16]
  assign _T_240 = {_T_228,_T_227}; // @[rvmemarb.scala 319:45:@4016.16]
  assign _T_241 = {_T_240,_T_221}; // @[rvmemarb.scala 319:45:@4017.16]
  assign _T_242 = 1'h0 == io_dm_port_req_mfunc; // @[Conditional.scala 37:30:@4023.10]
  assign _GEN_34 = io_dm_port_req_mfunc ? 1'h0 : _T_242; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_56 = io_dm_port_req_valid ? _GEN_34 : io_inst_port_req_valid; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_79 = reg_dmvld ? 1'h0 : 1'h1; // @[rvmemarb.scala 495:44:@4180.16]
  assign _GEN_81 = reg_rabusy ? 1'h0 : _GEN_79; // @[rvmemarb.scala 472:42:@4158.14]
  assign _GEN_98 = _T_242 ? _GEN_81 : 1'h0; // @[Conditional.scala 39:67:@4155.12]
  assign _GEN_115 = io_dm_port_req_mfunc ? 1'h0 : _GEN_98; // @[Conditional.scala 40:58:@4056.10]
  assign _GEN_131 = io_dm_port_req_valid ? _GEN_115 : 1'h0; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_140 = reg_ipvld ? 1'h0 : 1'h1; // @[rvmemarb.scala 621:44:@4296.16]
  assign _GEN_142 = reg_rabusy ? 1'h0 : _GEN_140; // @[rvmemarb.scala 598:42:@4274.14]
  assign _GEN_163 = io_inst_port_req_valid ? _GEN_142 : 1'h0; // @[rvmemarb.scala 588:42:@4270.10]
  assign _T_564 = 1'h0 == io_data_port_req_mfunc; // @[Conditional.scala 37:30:@4453.16]
  assign _GEN_188 = reg_dpvld ? 1'h0 : 1'h1; // @[rvmemarb.scala 823:44:@4479.20]
  assign _GEN_190 = reg_rabusy ? 1'h0 : _GEN_188; // @[rvmemarb.scala 800:42:@4457.18]
  assign _GEN_204 = _T_564 ? _GEN_190 : 1'h0; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_226 = io_data_port_req_mfunc ? 1'h0 : _GEN_204; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_244 = io_data_port_req_valid ? _GEN_226 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_262 = _T_467 ? _GEN_244 : 1'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_269 = _T_442 ? _GEN_163 : _GEN_262; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_296 = _T_252 ? _GEN_131 : _GEN_269; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_318 = _T_147 ? _GEN_56 : _GEN_296; // @[Conditional.scala 40:58:@3922.4]
  assign raen = reset ? 1'h0 : _GEN_318; // @[rvmemarb.scala 953:26:@4584.4]
  assign _T_245 = raen & io_ext_mem_rardy; // @[rvmemarb.scala 333:34:@4028.12]
  assign _GEN_20 = _T_245 ? 1'h1 : reg_rabusy; // @[rvmemarb.scala 333:42:@4029.12]
  assign _GEN_21 = _T_242 ? io_dm_port_req_addr : 32'h0; // @[Conditional.scala 39:67:@4024.10]
  assign _GEN_24 = _T_242 ? _GEN_20 : reg_rabusy; // @[Conditional.scala 39:67:@4024.10]
  assign _GEN_25 = io_dm_port_req_mfunc ? io_dm_port_req_addr : 32'h0; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_26 = io_dm_port_req_mfunc ? _GEN_13 : 1'h0; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_29 = io_dm_port_req_mfunc ? _GEN_11 : reg_wabusy; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_30 = io_dm_port_req_mfunc ? _GEN_12 : reg_wdbusy; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_31 = io_dm_port_req_mfunc ? _T_241 : 32'h0; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_32 = io_dm_port_req_mfunc ? 4'hf : 4'h0; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_33 = io_dm_port_req_mfunc ? 32'h0 : _GEN_21; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_36 = io_dm_port_req_mfunc ? reg_rabusy : _GEN_24; // @[Conditional.scala 40:58:@3925.8]
  assign _GEN_42 = io_inst_port_req_valid ? io_inst_port_req_addr : 32'h0; // @[rvmemarb.scala 341:47:@4036.8]
  assign _GEN_45 = io_inst_port_req_valid ? _GEN_20 : reg_rabusy; // @[rvmemarb.scala 341:47:@4036.8]
  assign _GEN_46 = io_inst_port_req_valid ? 2'h2 : reg_stat; // @[rvmemarb.scala 341:47:@4036.8]
  assign _GEN_47 = io_dm_port_req_valid ? _GEN_25 : 32'h0; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_48 = io_dm_port_req_valid ? _GEN_26 : 1'h0; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_51 = io_dm_port_req_valid ? _GEN_29 : reg_wabusy; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_52 = io_dm_port_req_valid ? _GEN_30 : reg_wdbusy; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_53 = io_dm_port_req_valid ? _GEN_31 : 32'h0; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_54 = io_dm_port_req_valid ? _GEN_32 : 4'h0; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_55 = io_dm_port_req_valid ? _GEN_33 : _GEN_42; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_58 = io_dm_port_req_valid ? _GEN_36 : _GEN_45; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_59 = io_dm_port_req_valid ? 2'h1 : _GEN_46; // @[rvmemarb.scala 225:40:@3923.6]
  assign _GEN_71 = io_ext_mem_rdrdy ? 1'h0 : reg_rabusy; // @[rvmemarb.scala 476:45:@4162.18]
  assign _GEN_72 = io_ext_mem_rdrdy ? 1'h0 : reg_rdbusy; // @[rvmemarb.scala 476:45:@4162.18]
  assign _GEN_74 = io_ext_mem_rdrdy ? 1'h0 : 1'h1; // @[rvmemarb.scala 486:45:@4171.18]
  assign _GEN_76 = reg_rdbusy ? _GEN_72 : _GEN_74; // @[rvmemarb.scala 475:46:@4161.16]
  assign _GEN_78 = reg_rdbusy ? 1'h0 : 1'h1; // @[rvmemarb.scala 475:46:@4161.16]
  assign _GEN_82 = reg_rabusy ? _GEN_78 : 1'h0; // @[rvmemarb.scala 472:42:@4158.14]
  assign _GEN_83 = reg_rabusy ? _GEN_71 : _GEN_20; // @[rvmemarb.scala 472:42:@4158.14]
  assign _GEN_84 = reg_rabusy ? _GEN_76 : reg_rdbusy; // @[rvmemarb.scala 472:42:@4158.14]
  assign _T_373 = io_ext_mem_rdata[7:0]; // @[rvmemarb.scala 514:88:@4193.18]
  assign _T_374 = {24'h0,_T_373}; // @[Cat.scala 30:58:@4194.18]
  assign _T_381 = io_ext_mem_rdata[15:8]; // @[rvmemarb.scala 515:88:@4196.18]
  assign _T_382 = {24'h0,_T_381}; // @[Cat.scala 30:58:@4197.18]
  assign _T_389 = io_ext_mem_rdata[23:16]; // @[rvmemarb.scala 516:88:@4199.18]
  assign _T_390 = {24'h0,_T_389}; // @[Cat.scala 30:58:@4200.18]
  assign _T_397 = io_ext_mem_rdata[31:24]; // @[rvmemarb.scala 517:88:@4202.18]
  assign _T_398 = {24'h0,_T_397}; // @[Cat.scala 30:58:@4203.18]
  assign _T_419 = {16'h0,_T_381}; // @[Cat.scala 30:58:@4222.20]
  assign _T_420 = {_T_419,_T_373}; // @[Cat.scala 30:58:@4223.20]
  assign _T_429 = {16'h0,_T_397}; // @[Cat.scala 30:58:@4227.20]
  assign _T_430 = {_T_429,_T_389}; // @[Cat.scala 30:58:@4228.20]
  assign _GEN_92 = io_ext_mem_rdrdy ? io_ext_mem_rdata : reg_dmdata; // @[rvmemarb.scala 505:37:@4189.14]
  assign _T_439 = io_dm_port_req_valid == 1'h0; // @[rvmemarb.scala 551:34:@4244.16]
  assign _GEN_94 = io_inst_port_req_valid ? 2'h2 : 2'h0; // @[rvmemarb.scala 552:62:@4246.18]
  assign _GEN_95 = _T_439 ? _GEN_94 : reg_stat; // @[rvmemarb.scala 551:57:@4245.16]
  assign _GEN_96 = reg_dmvld ? _GEN_95 : reg_stat; // @[rvmemarb.scala 546:40:@4243.14]
  assign _GEN_99 = _T_242 ? _GEN_82 : 1'h0; // @[Conditional.scala 39:67:@4155.12]
  assign _GEN_100 = _T_242 ? _GEN_83 : reg_rabusy; // @[Conditional.scala 39:67:@4155.12]
  assign _GEN_101 = _T_242 ? _GEN_84 : reg_rdbusy; // @[Conditional.scala 39:67:@4155.12]
  assign _GEN_103 = _T_242 ? _GEN_92 : reg_dmdata; // @[Conditional.scala 39:67:@4155.12]
  assign _GEN_104 = _T_242 ? io_ext_mem_rdrdy : 1'h0; // @[Conditional.scala 39:67:@4155.12]
  assign _GEN_105 = _T_242 ? _GEN_96 : reg_stat; // @[Conditional.scala 39:67:@4155.12]
  assign _GEN_107 = io_dm_port_req_mfunc ? _GEN_13 : 1'h1; // @[Conditional.scala 40:58:@4056.10]
  assign _GEN_116 = io_dm_port_req_mfunc ? 1'h0 : _GEN_99; // @[Conditional.scala 40:58:@4056.10]
  assign _GEN_117 = io_dm_port_req_mfunc ? reg_rabusy : _GEN_100; // @[Conditional.scala 40:58:@4056.10]
  assign _GEN_118 = io_dm_port_req_mfunc ? reg_rdbusy : _GEN_101; // @[Conditional.scala 40:58:@4056.10]
  assign _GEN_119 = io_dm_port_req_mfunc ? reg_dmdata : _GEN_103; // @[Conditional.scala 40:58:@4056.10]
  assign _GEN_120 = io_dm_port_req_mfunc ? 1'h0 : _GEN_104; // @[Conditional.scala 40:58:@4056.10]
  assign _GEN_121 = io_dm_port_req_mfunc ? reg_stat : _GEN_105; // @[Conditional.scala 40:58:@4056.10]
  assign _GEN_122 = io_dm_port_req_valid ? _GEN_107 : 1'h0; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_126 = io_dm_port_req_valid ? _GEN_29 : 1'h0; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_127 = io_dm_port_req_valid ? _GEN_30 : 1'h0; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_130 = io_dm_port_req_valid ? _GEN_33 : 32'h0; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_132 = io_dm_port_req_valid ? _GEN_116 : 1'h0; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_133 = io_dm_port_req_valid ? _GEN_117 : reg_rabusy; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_134 = io_dm_port_req_valid ? _GEN_118 : reg_rdbusy; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_135 = io_dm_port_req_valid ? _GEN_119 : reg_dmdata; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_136 = io_dm_port_req_valid ? _GEN_120 : 1'h0; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_137 = io_dm_port_req_valid ? _GEN_121 : _GEN_94; // @[rvmemarb.scala 361:40:@4053.8]
  assign _GEN_144 = reg_rabusy ? io_ext_mem_rdrdy : 1'h0; // @[rvmemarb.scala 598:42:@4274.14]
  assign _GEN_145 = io_ext_mem_rdrdy ? io_ext_mem_rdata : reg_ipdata; // @[rvmemarb.scala 632:37:@4305.14]
  assign _T_463 = io_inst_port_req_valid == 1'h0; // @[rvmemarb.scala 650:39:@4320.20]
  assign _GEN_146 = _T_463 ? 2'h0 : reg_stat; // @[rvmemarb.scala 650:64:@4321.20]
  assign _GEN_147 = io_dm_port_req_valid ? 2'h1 : _GEN_146; // @[rvmemarb.scala 647:61:@4316.18]
  assign _GEN_148 = io_data_port_req_valid ? 2'h3 : _GEN_147; // @[rvmemarb.scala 643:58:@4311.16]
  assign _GEN_149 = io_data_port_req_valid ? 1'h1 : io_ext_mem_rdrdy; // @[rvmemarb.scala 643:58:@4311.16]
  assign _GEN_150 = reg_ipvld ? 1'h0 : _GEN_84; // @[rvmemarb.scala 638:40:@4309.14]
  assign _GEN_151 = reg_ipvld ? _GEN_148 : reg_stat; // @[rvmemarb.scala 638:40:@4309.14]
  assign _GEN_152 = reg_ipvld ? _GEN_149 : io_ext_mem_rdrdy; // @[rvmemarb.scala 638:40:@4309.14]
  assign _GEN_164 = io_inst_port_req_valid ? _GEN_82 : 1'h0; // @[rvmemarb.scala 588:42:@4270.10]
  assign _GEN_165 = io_inst_port_req_valid ? _GEN_83 : reg_rabusy; // @[rvmemarb.scala 588:42:@4270.10]
  assign _GEN_166 = io_inst_port_req_valid ? _GEN_150 : reg_rdbusy; // @[rvmemarb.scala 588:42:@4270.10]
  assign _GEN_168 = io_inst_port_req_valid ? _GEN_152 : 1'h0; // @[rvmemarb.scala 588:42:@4270.10]
  assign _GEN_169 = io_inst_port_req_valid ? _GEN_145 : 32'h13; // @[rvmemarb.scala 588:42:@4270.10]
  assign _GEN_170 = io_inst_port_req_valid ? _GEN_151 : 2'h0; // @[rvmemarb.scala 588:42:@4270.10]
  assign _GEN_171 = io_inst_port_req_valid ? reg_wabusy : 1'h0; // @[rvmemarb.scala 588:42:@4270.10]
  assign _GEN_172 = io_inst_port_req_valid ? reg_wdbusy : 1'h0; // @[rvmemarb.scala 588:42:@4270.10]
  assign _T_470 = io_data_port_req_addr[1:0]; // @[rvmemarb.scala 684:48:@4342.16]
  assign _T_484 = 2'h1 == io_data_port_req_mtype; // @[Conditional.scala 37:30:@4371.16]
  assign _T_485 = io_data_port_req_data[7:0]; // @[rvmemarb.scala 721:41:@4373.18]
  assign _T_507 = 2'h3 == _T_470; // @[Mux.scala 46:19:@4382.18]
  assign _T_508 = _T_507 ? 4'h8 : 4'h0; // @[Mux.scala 46:16:@4383.18]
  assign _T_509 = 2'h2 == _T_470; // @[Mux.scala 46:19:@4384.18]
  assign _T_510 = _T_509 ? 4'h4 : _T_508; // @[Mux.scala 46:16:@4385.18]
  assign _T_511 = 2'h1 == _T_470; // @[Mux.scala 46:19:@4386.18]
  assign _T_512 = _T_511 ? 4'h2 : _T_510; // @[Mux.scala 46:16:@4387.18]
  assign _T_513 = 2'h0 == _T_470; // @[Mux.scala 46:19:@4388.18]
  assign _T_514 = _T_513 ? 4'h1 : _T_512; // @[Mux.scala 46:16:@4389.18]
  assign _T_515 = {_T_485,_T_485}; // @[rvmemarb.scala 737:45:@4390.18]
  assign _T_517 = {_T_515,_T_515}; // @[rvmemarb.scala 737:45:@4392.18]
  assign _T_518 = 2'h2 == io_data_port_req_mtype; // @[Conditional.scala 37:30:@4397.18]
  assign _T_520 = io_data_port_req_data[15:8]; // @[rvmemarb.scala 744:41:@4400.20]
  assign _T_532 = _T_470[1]; // @[rvmemarb.scala 749:40:@4408.20]
  assign _T_539 = _T_532 ? 4'hc : 4'h0; // @[Mux.scala 46:16:@4410.20]
  assign _T_540 = 1'h0 == _T_532; // @[Mux.scala 46:19:@4411.20]
  assign _T_541 = _T_540 ? 4'h3 : _T_539; // @[Mux.scala 46:16:@4412.20]
  assign _T_542 = {_T_520,_T_485}; // @[rvmemarb.scala 757:45:@4413.20]
  assign _T_544 = {_T_542,_T_542}; // @[rvmemarb.scala 757:45:@4415.20]
  assign _T_545 = 2'h3 == io_data_port_req_mtype; // @[Conditional.scala 37:30:@4420.20]
  assign _T_548 = io_data_port_req_data[23:16]; // @[rvmemarb.scala 765:41:@4424.22]
  assign _T_549 = io_data_port_req_data[31:24]; // @[rvmemarb.scala 766:41:@4425.22]
  assign _T_561 = {_T_549,_T_548}; // @[rvmemarb.scala 770:45:@4432.22]
  assign _T_562 = {_T_561,_T_542}; // @[rvmemarb.scala 770:45:@4433.22]
  assign _GEN_178 = _T_545 ? _T_562 : 32'h0; // @[Conditional.scala 39:67:@4421.20]
  assign _GEN_179 = _T_545 ? 4'hf : 4'h0; // @[Conditional.scala 39:67:@4421.20]
  assign _GEN_180 = _T_518 ? _T_544 : _GEN_178; // @[Conditional.scala 39:67:@4398.18]
  assign _GEN_181 = _T_518 ? _T_541 : _GEN_179; // @[Conditional.scala 39:67:@4398.18]
  assign _GEN_182 = _T_484 ? _T_517 : _GEN_180; // @[Conditional.scala 40:58:@4372.16]
  assign _GEN_183 = _T_484 ? _T_514 : _GEN_181; // @[Conditional.scala 40:58:@4372.16]
  assign _GEN_184 = io_dm_port_req_valid ? 2'h1 : _GEN_94; // @[rvmemarb.scala 783:56:@4440.18]
  assign _GEN_185 = io_ext_mem_wbvld ? 1'h0 : 1'h1; // @[rvmemarb.scala 780:37:@4437.16]
  assign _GEN_186 = io_ext_mem_wbvld ? 32'h13 : reg_ipdata; // @[rvmemarb.scala 780:37:@4437.16]
  assign _GEN_187 = io_ext_mem_wbvld ? _GEN_184 : reg_stat; // @[rvmemarb.scala 780:37:@4437.16]
  assign _T_616 = _T_507 ? _T_398 : 32'h0; // @[Mux.scala 46:16:@4504.22]
  assign _T_618 = _T_509 ? _T_390 : _T_616; // @[Mux.scala 46:16:@4506.22]
  assign _T_620 = _T_511 ? _T_382 : _T_618; // @[Mux.scala 46:16:@4508.22]
  assign _T_622 = _T_513 ? _T_374 : _T_620; // @[Mux.scala 46:16:@4510.22]
  assign _T_648 = _T_532 ? _T_430 : 32'h0; // @[Mux.scala 46:16:@4529.24]
  assign _T_650 = _T_540 ? _T_420 : _T_648; // @[Mux.scala 46:16:@4531.24]
  assign _GEN_192 = _T_545 ? io_ext_mem_rdata : reg_dpdata; // @[Conditional.scala 39:67:@4537.24]
  assign _GEN_194 = _T_518 ? _T_650 : _GEN_192; // @[Conditional.scala 39:67:@4516.22]
  assign _GEN_195 = _T_518 ? 1'h1 : _T_545; // @[Conditional.scala 39:67:@4516.22]
  assign _GEN_196 = _T_484 ? _T_622 : _GEN_194; // @[Conditional.scala 40:58:@4490.20]
  assign _GEN_197 = _T_484 ? 1'h1 : _GEN_195; // @[Conditional.scala 40:58:@4490.20]
  assign _GEN_198 = io_ext_mem_rdrdy ? _GEN_196 : reg_dpdata; // @[rvmemarb.scala 834:37:@4488.18]
  assign _GEN_199 = io_ext_mem_rdrdy ? _GEN_197 : 1'h0; // @[rvmemarb.scala 834:37:@4488.18]
  assign _GEN_200 = reg_dpvld ? 1'h0 : _GEN_84; // @[rvmemarb.scala 876:40:@4542.18]
  assign _GEN_201 = reg_dpvld ? 32'h13 : reg_ipdata; // @[rvmemarb.scala 876:40:@4542.18]
  assign _GEN_202 = reg_dpvld ? _GEN_184 : reg_stat; // @[rvmemarb.scala 876:40:@4542.18]
  assign _GEN_203 = _T_564 ? io_data_port_req_addr : 32'h0; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_205 = _T_564 ? _GEN_82 : 1'h0; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_206 = _T_564 ? _GEN_83 : reg_rabusy; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_207 = _T_564 ? _GEN_200 : reg_rdbusy; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_208 = _T_564 ? _GEN_144 : 1'h0; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_209 = _T_564 ? _GEN_198 : reg_dpdata; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_210 = _T_564 ? _GEN_199 : 1'h0; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_211 = _T_564 ? _GEN_188 : 1'h1; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_212 = _T_564 ? _GEN_201 : reg_ipdata; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_213 = _T_564 ? _GEN_202 : reg_stat; // @[Conditional.scala 39:67:@4454.16]
  assign _GEN_214 = io_data_port_req_mfunc ? io_data_port_req_addr : 32'h0; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_215 = io_data_port_req_mfunc ? _GEN_13 : _GEN_208; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_218 = io_data_port_req_mfunc ? _GEN_11 : reg_wabusy; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_219 = io_data_port_req_mfunc ? _GEN_12 : reg_wdbusy; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_220 = io_data_port_req_mfunc ? _GEN_182 : 32'h0; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_221 = io_data_port_req_mfunc ? _GEN_183 : 4'h0; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_222 = io_data_port_req_mfunc ? _GEN_185 : _GEN_211; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_223 = io_data_port_req_mfunc ? _GEN_186 : _GEN_212; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_224 = io_data_port_req_mfunc ? _GEN_187 : _GEN_213; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_225 = io_data_port_req_mfunc ? 32'h0 : _GEN_203; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_227 = io_data_port_req_mfunc ? 1'h0 : _GEN_205; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_228 = io_data_port_req_mfunc ? reg_rabusy : _GEN_206; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_229 = io_data_port_req_mfunc ? reg_rdbusy : _GEN_207; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_230 = io_data_port_req_mfunc ? reg_dpdata : _GEN_209; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_231 = io_data_port_req_mfunc ? 1'h0 : _GEN_210; // @[Conditional.scala 40:58:@4341.14]
  assign _GEN_232 = io_data_port_req_valid ? _GEN_214 : 32'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_233 = io_data_port_req_valid ? _GEN_215 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_236 = io_data_port_req_valid ? _GEN_218 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_237 = io_data_port_req_valid ? _GEN_219 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_238 = io_data_port_req_valid ? _GEN_220 : 32'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_239 = io_data_port_req_valid ? _GEN_221 : 4'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_240 = io_data_port_req_valid ? _GEN_222 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_241 = io_data_port_req_valid ? _GEN_223 : 32'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_242 = io_data_port_req_valid ? _GEN_224 : 2'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_243 = io_data_port_req_valid ? _GEN_225 : 32'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_245 = io_data_port_req_valid ? _GEN_227 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_246 = io_data_port_req_valid ? _GEN_228 : reg_rabusy; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_247 = io_data_port_req_valid ? _GEN_229 : reg_rdbusy; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_248 = io_data_port_req_valid ? _GEN_230 : reg_dpdata; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_249 = io_data_port_req_valid ? _GEN_231 : 1'h0; // @[rvmemarb.scala 677:42:@4339.12]
  assign _GEN_250 = _T_467 ? _GEN_240 : 1'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_251 = _T_467 ? _GEN_232 : 32'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_252 = _T_467 ? _GEN_233 : 1'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_255 = _T_467 ? _GEN_236 : reg_wabusy; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_256 = _T_467 ? _GEN_237 : reg_wdbusy; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_257 = _T_467 ? _GEN_238 : 32'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_258 = _T_467 ? _GEN_239 : 4'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_259 = _T_467 ? _GEN_241 : reg_ipdata; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_260 = _T_467 ? _GEN_242 : reg_stat; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_261 = _T_467 ? _GEN_243 : 32'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_263 = _T_467 ? _GEN_245 : 1'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_264 = _T_467 ? _GEN_246 : reg_rabusy; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_265 = _T_467 ? _GEN_247 : reg_rdbusy; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_266 = _T_467 ? _GEN_248 : reg_dpdata; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_267 = _T_467 ? _GEN_249 : 1'h0; // @[Conditional.scala 39:67:@4337.10]
  assign _GEN_268 = _T_442 ? _GEN_42 : _GEN_261; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_270 = _T_442 ? _GEN_164 : _GEN_263; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_271 = _T_442 ? _GEN_165 : _GEN_264; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_272 = _T_442 ? _GEN_166 : _GEN_265; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_274 = _T_442 ? _GEN_168 : _GEN_250; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_275 = _T_442 ? _GEN_169 : _GEN_259; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_276 = _T_442 ? _GEN_170 : _GEN_260; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_277 = _T_442 ? _GEN_171 : _GEN_255; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_278 = _T_442 ? _GEN_172 : _GEN_256; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_279 = _T_442 ? 32'h0 : _GEN_251; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_280 = _T_442 ? 1'h0 : _GEN_252; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_283 = _T_442 ? 32'h0 : _GEN_257; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_284 = _T_442 ? 4'h0 : _GEN_258; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_285 = _T_442 ? reg_dpdata : _GEN_266; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_286 = _T_442 ? 1'h0 : _GEN_267; // @[Conditional.scala 39:67:@4269.8]
  assign _GEN_287 = _T_252 ? _GEN_122 : 1'h0; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_288 = _T_252 ? _GEN_47 : _GEN_279; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_291 = _T_252 ? _GEN_126 : _GEN_277; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_292 = _T_252 ? _GEN_127 : _GEN_278; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_293 = _T_252 ? _GEN_53 : _GEN_283; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_294 = _T_252 ? _GEN_54 : _GEN_284; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_295 = _T_252 ? _GEN_130 : _GEN_268; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_297 = _T_252 ? _GEN_132 : _GEN_270; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_298 = _T_252 ? _GEN_133 : _GEN_271; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_299 = _T_252 ? _GEN_134 : _GEN_272; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_300 = _T_252 ? _GEN_135 : reg_dmdata; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_301 = _T_252 ? _GEN_136 : 1'h0; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_302 = _T_252 ? _GEN_137 : _GEN_276; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_304 = _T_252 ? 1'h0 : _GEN_274; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_305 = _T_252 ? reg_ipdata : _GEN_275; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_306 = _T_252 ? 1'h0 : _GEN_280; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_307 = _T_252 ? reg_dpdata : _GEN_285; // @[Conditional.scala 39:67:@4052.6]
  assign _GEN_308 = _T_252 ? 1'h0 : _GEN_286; // @[Conditional.scala 39:67:@4052.6]
  assign waddr = _T_147 ? _GEN_47 : _GEN_288; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_310 = _T_147 ? _GEN_48 : _GEN_287; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_313 = _T_147 ? _GEN_51 : _GEN_291; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_314 = _T_147 ? _GEN_52 : _GEN_292; // @[Conditional.scala 40:58:@3922.4]
  assign wdata = _T_147 ? _GEN_53 : _GEN_293; // @[Conditional.scala 40:58:@3922.4]
  assign wmask = _T_147 ? _GEN_54 : _GEN_294; // @[Conditional.scala 40:58:@3922.4]
  assign raddr = _T_147 ? _GEN_55 : _GEN_295; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_319 = _T_147 ? 1'h0 : _GEN_297; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_320 = _T_147 ? _GEN_58 : _GEN_298; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_321 = _T_147 ? _GEN_59 : _GEN_302; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_322 = _T_147 ? reg_rdbusy : _GEN_299; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_323 = _T_147 ? reg_dmdata : _GEN_300; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_324 = _T_147 ? 1'h0 : _GEN_301; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_326 = _T_147 ? 1'h0 : _GEN_304; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_327 = _T_147 ? reg_ipdata : _GEN_305; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_328 = _T_147 ? 1'h0 : _GEN_306; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_329 = _T_147 ? reg_dpdata : _GEN_307; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_330 = _T_147 ? 1'h0 : _GEN_308; // @[Conditional.scala 40:58:@3922.4]
  assign _GEN_331 = reset ? 2'h0 : _GEN_321; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_332 = reset ? 1'h0 : _GEN_313; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_333 = reset ? 1'h0 : _GEN_314; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_334 = reset ? 1'h0 : _GEN_320; // @[rvmemarb.scala 953:26:@4584.4]
  assign rden = reset ? 1'h0 : _GEN_319; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_340 = reset ? 1'h0 : _GEN_328; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_341 = reset ? 1'h0 : _GEN_310; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_342 = reset ? 1'h0 : reg_ipvld; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_343 = reset ? 1'h0 : reg_dpvld; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_344 = reset ? 1'h0 : reg_dmvld; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_345 = reset ? 32'h0 : _GEN_323; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_346 = reset ? 1'h0 : _GEN_324; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_347 = reset ? 32'h0 : _GEN_327; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_348 = reset ? 1'h0 : _GEN_326; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_349 = reset ? 32'h0 : _GEN_329; // @[rvmemarb.scala 953:26:@4584.4]
  assign _GEN_350 = reset ? 1'h0 : _GEN_330; // @[rvmemarb.scala 953:26:@4584.4]
  assign io_inst_port_resp_data = reg_ipdata;
  assign io_inst_port_resp_valid = _GEN_342;
  assign io_data_port_req_ready = _GEN_340;
  assign io_data_port_resp_data = reg_dpdata;
  assign io_data_port_resp_valid = _GEN_343;
  assign io_dm_port_req_ready = _GEN_341;
  assign io_dm_port_resp_data = reg_dmdata;
  assign io_dm_port_resp_valid = _GEN_344;
  assign io_ext_mem_waen = waen;
  assign io_ext_mem_wden = wden;
  assign io_ext_mem_waddr = waddr;
  assign io_ext_mem_wdata = wdata;
  assign io_ext_mem_wmask = wmask;
  assign io_ext_mem_raen = raen;
  assign io_ext_mem_rden = rden;
  assign io_ext_mem_raddr = raddr;
  assign io_ext_mem_clock = clock;
  assign io_ext_mem_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  reg_stat = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  reg_wabusy = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  reg_wdbusy = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  reg_rabusy = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  reg_rdbusy = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  reg_dmdata = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  reg_dmvld = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  reg_ipdata = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  reg_ipvld = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  reg_dpdata = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  reg_dpvld = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_stat <= 2'h0;
    end else begin
      if (_T_147) begin
        if (io_dm_port_req_valid) begin
          reg_stat <= 2'h1;
        end else begin
          if (io_inst_port_req_valid) begin
            reg_stat <= 2'h2;
          end
        end
      end else begin
        if (_T_252) begin
          if (io_dm_port_req_valid) begin
            if (!(io_dm_port_req_mfunc)) begin
              if (_T_242) begin
                if (reg_dmvld) begin
                  if (_T_439) begin
                    if (io_inst_port_req_valid) begin
                      reg_stat <= 2'h2;
                    end else begin
                      reg_stat <= 2'h0;
                    end
                  end
                end
              end
            end
          end else begin
            if (io_inst_port_req_valid) begin
              reg_stat <= 2'h2;
            end else begin
              reg_stat <= 2'h0;
            end
          end
        end else begin
          if (_T_442) begin
            if (io_inst_port_req_valid) begin
              if (reg_ipvld) begin
                if (io_data_port_req_valid) begin
                  reg_stat <= 2'h3;
                end else begin
                  if (io_dm_port_req_valid) begin
                    reg_stat <= 2'h1;
                  end else begin
                    if (_T_463) begin
                      reg_stat <= 2'h0;
                    end
                  end
                end
              end
            end else begin
              reg_stat <= 2'h0;
            end
          end else begin
            if (_T_467) begin
              if (io_data_port_req_valid) begin
                if (io_data_port_req_mfunc) begin
                  if (io_ext_mem_wbvld) begin
                    if (io_dm_port_req_valid) begin
                      reg_stat <= 2'h1;
                    end else begin
                      if (io_inst_port_req_valid) begin
                        reg_stat <= 2'h2;
                      end else begin
                        reg_stat <= 2'h0;
                      end
                    end
                  end
                end else begin
                  if (_T_564) begin
                    if (reg_dpvld) begin
                      if (io_dm_port_req_valid) begin
                        reg_stat <= 2'h1;
                      end else begin
                        if (io_inst_port_req_valid) begin
                          reg_stat <= 2'h2;
                        end else begin
                          reg_stat <= 2'h0;
                        end
                      end
                    end
                  end
                end
              end else begin
                reg_stat <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_wabusy <= 1'h0;
    end else begin
      if (_T_147) begin
        if (io_dm_port_req_valid) begin
          if (io_dm_port_req_mfunc) begin
            if (reg_wabusy) begin
              if (reg_wdbusy) begin
                if (io_ext_mem_wbvld) begin
                  reg_wabusy <= 1'h0;
                end
              end
            end else begin
              if (_T_161) begin
                reg_wabusy <= 1'h1;
              end
            end
          end
        end
      end else begin
        if (_T_252) begin
          if (io_dm_port_req_valid) begin
            if (io_dm_port_req_mfunc) begin
              if (reg_wabusy) begin
                if (reg_wdbusy) begin
                  if (io_ext_mem_wbvld) begin
                    reg_wabusy <= 1'h0;
                  end
                end
              end else begin
                if (_T_161) begin
                  reg_wabusy <= 1'h1;
                end
              end
            end
          end else begin
            reg_wabusy <= 1'h0;
          end
        end else begin
          if (_T_442) begin
            if (!(io_inst_port_req_valid)) begin
              reg_wabusy <= 1'h0;
            end
          end else begin
            if (_T_467) begin
              if (io_data_port_req_valid) begin
                if (io_data_port_req_mfunc) begin
                  if (reg_wabusy) begin
                    if (reg_wdbusy) begin
                      if (io_ext_mem_wbvld) begin
                        reg_wabusy <= 1'h0;
                      end
                    end
                  end else begin
                    if (_T_161) begin
                      reg_wabusy <= 1'h1;
                    end
                  end
                end
              end else begin
                reg_wabusy <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_wdbusy <= 1'h0;
    end else begin
      if (_T_147) begin
        if (io_dm_port_req_valid) begin
          if (io_dm_port_req_mfunc) begin
            if (reg_wabusy) begin
              if (reg_wdbusy) begin
                if (io_ext_mem_wbvld) begin
                  reg_wdbusy <= 1'h0;
                end
              end else begin
                if (_T_157) begin
                  reg_wdbusy <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_252) begin
          if (io_dm_port_req_valid) begin
            if (io_dm_port_req_mfunc) begin
              if (reg_wabusy) begin
                if (reg_wdbusy) begin
                  if (io_ext_mem_wbvld) begin
                    reg_wdbusy <= 1'h0;
                  end
                end else begin
                  if (_T_157) begin
                    reg_wdbusy <= 1'h1;
                  end
                end
              end
            end
          end else begin
            reg_wdbusy <= 1'h0;
          end
        end else begin
          if (_T_442) begin
            if (!(io_inst_port_req_valid)) begin
              reg_wdbusy <= 1'h0;
            end
          end else begin
            if (_T_467) begin
              if (io_data_port_req_valid) begin
                if (io_data_port_req_mfunc) begin
                  if (reg_wabusy) begin
                    if (reg_wdbusy) begin
                      if (io_ext_mem_wbvld) begin
                        reg_wdbusy <= 1'h0;
                      end
                    end else begin
                      if (_T_157) begin
                        reg_wdbusy <= 1'h1;
                      end
                    end
                  end
                end
              end else begin
                reg_wdbusy <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_rabusy <= 1'h0;
    end else begin
      if (_T_147) begin
        if (io_dm_port_req_valid) begin
          if (!(io_dm_port_req_mfunc)) begin
            if (_T_242) begin
              if (_T_245) begin
                reg_rabusy <= 1'h1;
              end
            end
          end
        end else begin
          if (io_inst_port_req_valid) begin
            if (_T_245) begin
              reg_rabusy <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_252) begin
          if (io_dm_port_req_valid) begin
            if (!(io_dm_port_req_mfunc)) begin
              if (_T_242) begin
                if (reg_rabusy) begin
                  if (io_ext_mem_rdrdy) begin
                    reg_rabusy <= 1'h0;
                  end
                end else begin
                  if (_T_245) begin
                    reg_rabusy <= 1'h1;
                  end
                end
              end
            end
          end
        end else begin
          if (_T_442) begin
            if (io_inst_port_req_valid) begin
              if (reg_rabusy) begin
                if (io_ext_mem_rdrdy) begin
                  reg_rabusy <= 1'h0;
                end
              end else begin
                if (_T_245) begin
                  reg_rabusy <= 1'h1;
                end
              end
            end
          end else begin
            if (_T_467) begin
              if (io_data_port_req_valid) begin
                if (!(io_data_port_req_mfunc)) begin
                  if (_T_564) begin
                    if (reg_rabusy) begin
                      if (io_ext_mem_rdrdy) begin
                        reg_rabusy <= 1'h0;
                      end
                    end else begin
                      reg_rabusy <= _GEN_20;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (!(_T_147)) begin
      if (_T_252) begin
        if (io_dm_port_req_valid) begin
          if (!(io_dm_port_req_mfunc)) begin
            if (_T_242) begin
              if (reg_rabusy) begin
                if (reg_rdbusy) begin
                  if (io_ext_mem_rdrdy) begin
                    reg_rdbusy <= 1'h0;
                  end
                end else begin
                  if (io_ext_mem_rdrdy) begin
                    reg_rdbusy <= 1'h0;
                  end else begin
                    reg_rdbusy <= 1'h1;
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_442) begin
          if (io_inst_port_req_valid) begin
            if (reg_ipvld) begin
              reg_rdbusy <= 1'h0;
            end else begin
              if (reg_rabusy) begin
                if (reg_rdbusy) begin
                  if (io_ext_mem_rdrdy) begin
                    reg_rdbusy <= 1'h0;
                  end
                end else begin
                  if (io_ext_mem_rdrdy) begin
                    reg_rdbusy <= 1'h0;
                  end else begin
                    reg_rdbusy <= 1'h1;
                  end
                end
              end
            end
          end
        end else begin
          if (_T_467) begin
            if (io_data_port_req_valid) begin
              if (!(io_data_port_req_mfunc)) begin
                if (_T_564) begin
                  if (reg_dpvld) begin
                    reg_rdbusy <= 1'h0;
                  end else begin
                    if (reg_rabusy) begin
                      if (reg_rdbusy) begin
                        if (io_ext_mem_rdrdy) begin
                          reg_rdbusy <= 1'h0;
                        end
                      end else begin
                        if (io_ext_mem_rdrdy) begin
                          reg_rdbusy <= 1'h0;
                        end else begin
                          reg_rdbusy <= 1'h1;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dmdata <= 32'h0;
    end else begin
      if (!(_T_147)) begin
        if (_T_252) begin
          if (io_dm_port_req_valid) begin
            if (!(io_dm_port_req_mfunc)) begin
              if (_T_242) begin
                if (io_ext_mem_rdrdy) begin
                  reg_dmdata <= io_ext_mem_rdata;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dmvld <= 1'h0;
    end else begin
      if (_T_147) begin
        reg_dmvld <= 1'h0;
      end else begin
        if (_T_252) begin
          if (io_dm_port_req_valid) begin
            if (io_dm_port_req_mfunc) begin
              reg_dmvld <= 1'h0;
            end else begin
              if (_T_242) begin
                reg_dmvld <= io_ext_mem_rdrdy;
              end else begin
                reg_dmvld <= 1'h0;
              end
            end
          end else begin
            reg_dmvld <= 1'h0;
          end
        end else begin
          reg_dmvld <= 1'h0;
        end
      end
    end
    if (reset) begin
      reg_ipdata <= 32'h0;
    end else begin
      if (!(_T_147)) begin
        if (!(_T_252)) begin
          if (_T_442) begin
            if (io_inst_port_req_valid) begin
              if (io_ext_mem_rdrdy) begin
                reg_ipdata <= io_ext_mem_rdata;
              end
            end else begin
              reg_ipdata <= 32'h13;
            end
          end else begin
            if (_T_467) begin
              if (io_data_port_req_valid) begin
                if (io_data_port_req_mfunc) begin
                  if (io_ext_mem_wbvld) begin
                    reg_ipdata <= 32'h13;
                  end
                end else begin
                  if (_T_564) begin
                    if (reg_dpvld) begin
                      reg_ipdata <= 32'h13;
                    end
                  end
                end
              end else begin
                reg_ipdata <= 32'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_ipvld <= 1'h0;
    end else begin
      if (_T_147) begin
        reg_ipvld <= 1'h0;
      end else begin
        if (_T_252) begin
          reg_ipvld <= 1'h0;
        end else begin
          if (_T_442) begin
            if (io_inst_port_req_valid) begin
              if (reg_ipvld) begin
                if (io_data_port_req_valid) begin
                  reg_ipvld <= 1'h1;
                end else begin
                  reg_ipvld <= io_ext_mem_rdrdy;
                end
              end else begin
                reg_ipvld <= io_ext_mem_rdrdy;
              end
            end else begin
              reg_ipvld <= 1'h0;
            end
          end else begin
            if (_T_467) begin
              if (io_data_port_req_valid) begin
                if (io_data_port_req_mfunc) begin
                  if (io_ext_mem_wbvld) begin
                    reg_ipvld <= 1'h0;
                  end else begin
                    reg_ipvld <= 1'h1;
                  end
                end else begin
                  if (_T_564) begin
                    if (reg_dpvld) begin
                      reg_ipvld <= 1'h0;
                    end else begin
                      reg_ipvld <= 1'h1;
                    end
                  end else begin
                    reg_ipvld <= 1'h1;
                  end
                end
              end else begin
                reg_ipvld <= 1'h0;
              end
            end else begin
              reg_ipvld <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dpdata <= 32'h0;
    end else begin
      if (!(_T_147)) begin
        if (!(_T_252)) begin
          if (!(_T_442)) begin
            if (_T_467) begin
              if (io_data_port_req_valid) begin
                if (!(io_data_port_req_mfunc)) begin
                  if (_T_564) begin
                    if (io_ext_mem_rdrdy) begin
                      if (_T_484) begin
                        if (_T_513) begin
                          reg_dpdata <= _T_374;
                        end else begin
                          if (_T_511) begin
                            reg_dpdata <= _T_382;
                          end else begin
                            if (_T_509) begin
                              reg_dpdata <= _T_390;
                            end else begin
                              if (_T_507) begin
                                reg_dpdata <= _T_398;
                              end else begin
                                reg_dpdata <= 32'h0;
                              end
                            end
                          end
                        end
                      end else begin
                        if (_T_518) begin
                          if (_T_540) begin
                            reg_dpdata <= _T_420;
                          end else begin
                            if (_T_532) begin
                              reg_dpdata <= _T_430;
                            end else begin
                              reg_dpdata <= 32'h0;
                            end
                          end
                        end else begin
                          if (_T_545) begin
                            reg_dpdata <= io_ext_mem_rdata;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dpvld <= 1'h0;
    end else begin
      if (_T_147) begin
        reg_dpvld <= 1'h0;
      end else begin
        if (_T_252) begin
          reg_dpvld <= 1'h0;
        end else begin
          if (_T_442) begin
            reg_dpvld <= 1'h0;
          end else begin
            if (_T_467) begin
              if (io_data_port_req_valid) begin
                if (io_data_port_req_mfunc) begin
                  reg_dpvld <= 1'h0;
                end else begin
                  if (_T_564) begin
                    if (io_ext_mem_rdrdy) begin
                      if (_T_484) begin
                        reg_dpvld <= 1'h1;
                      end else begin
                        if (_T_518) begin
                          reg_dpvld <= 1'h1;
                        end else begin
                          reg_dpvld <= _T_545;
                        end
                      end
                    end else begin
                      reg_dpvld <= 1'h0;
                    end
                  end else begin
                    reg_dpvld <= 1'h0;
                  end
                end
              end else begin
                reg_dpvld <= 1'h0;
              end
            end else begin
              reg_dpvld <= 1'h0;
            end
          end
        end
      end
    end
  end
endmodule
module rvtile( // @[:@4608.2]
  input         clock, // @[:@4609.4]
  input         reset, // @[:@4610.4]
  input  [1:0]  io_dmi_req_bits_op, // @[:@4611.4]
  input  [6:0]  io_dmi_req_bits_addr, // @[:@4611.4]
  input  [31:0] io_dmi_req_bits_data, // @[:@4611.4]
  input         io_dmi_req_valid, // @[:@4611.4]
  output        io_dmi_req_ready, // @[:@4611.4]
  output [1:0]  io_dmi_resp_bits_resp, // @[:@4611.4]
  output [31:0] io_dmi_resp_bits_data, // @[:@4611.4]
  output        io_dmi_resp_valid, // @[:@4611.4]
  output        io_ext_mem_waen, // @[:@4611.4]
  output        io_ext_mem_wden, // @[:@4611.4]
  output [31:0] io_ext_mem_waddr, // @[:@4611.4]
  output [31:0] io_ext_mem_wdata, // @[:@4611.4]
  output [3:0]  io_ext_mem_wmask, // @[:@4611.4]
  input         io_ext_mem_wardy, // @[:@4611.4]
  input         io_ext_mem_wdrdy, // @[:@4611.4]
  input         io_ext_mem_wbvld, // @[:@4611.4]
  output        io_ext_mem_raen, // @[:@4611.4]
  output        io_ext_mem_rden, // @[:@4611.4]
  output [31:0] io_ext_mem_raddr, // @[:@4611.4]
  input  [31:0] io_ext_mem_rdata, // @[:@4611.4]
  input         io_ext_mem_rardy, // @[:@4611.4]
  input         io_ext_mem_rdrdy, // @[:@4611.4]
  output        io_ext_mem_clock, // @[:@4611.4]
  output        io_ext_mem_reset // @[:@4611.4]
);
  wire  dm_clock; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_reset; // @[rvtile.scala 29:20:@4613.4]
  wire [1:0] dm_io_dmi_req_bits_op; // @[rvtile.scala 29:20:@4613.4]
  wire [6:0] dm_io_dmi_req_bits_addr; // @[rvtile.scala 29:20:@4613.4]
  wire [31:0] dm_io_dmi_req_bits_data; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_dmi_req_valid; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_dmi_req_ready; // @[rvtile.scala 29:20:@4613.4]
  wire [1:0] dm_io_dmi_resp_bits_resp; // @[rvtile.scala 29:20:@4613.4]
  wire [31:0] dm_io_dmi_resp_bits_data; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_dmi_resp_valid; // @[rvtile.scala 29:20:@4613.4]
  wire [4:0] dm_io_ddpath_addr; // @[rvtile.scala 29:20:@4613.4]
  wire [31:0] dm_io_ddpath_wdata; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_ddpath_valid; // @[rvtile.scala 29:20:@4613.4]
  wire [31:0] dm_io_ddpath_rdata; // @[rvtile.scala 29:20:@4613.4]
  wire [31:0] dm_io_ddmem_req_addr; // @[rvtile.scala 29:20:@4613.4]
  wire [31:0] dm_io_ddmem_req_data; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_ddmem_req_mfunc; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_ddmem_req_valid; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_ddmem_req_ready; // @[rvtile.scala 29:20:@4613.4]
  wire [31:0] dm_io_ddmem_resp_data; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_ddmem_resp_valid; // @[rvtile.scala 29:20:@4613.4]
  wire  dm_io_rstcore; // @[rvtile.scala 29:20:@4613.4]
  wire  core_clock; // @[rvtile.scala 30:22:@4616.4]
  wire  core_reset; // @[rvtile.scala 30:22:@4616.4]
  wire [31:0] core_io_imem_req_addr; // @[rvtile.scala 30:22:@4616.4]
  wire  core_io_imem_req_valid; // @[rvtile.scala 30:22:@4616.4]
  wire [31:0] core_io_imem_resp_data; // @[rvtile.scala 30:22:@4616.4]
  wire  core_io_imem_resp_valid; // @[rvtile.scala 30:22:@4616.4]
  wire [31:0] core_io_dmem_req_addr; // @[rvtile.scala 30:22:@4616.4]
  wire [31:0] core_io_dmem_req_data; // @[rvtile.scala 30:22:@4616.4]
  wire  core_io_dmem_req_mfunc; // @[rvtile.scala 30:22:@4616.4]
  wire [1:0] core_io_dmem_req_mtype; // @[rvtile.scala 30:22:@4616.4]
  wire  core_io_dmem_req_valid; // @[rvtile.scala 30:22:@4616.4]
  wire  core_io_dmem_req_ready; // @[rvtile.scala 30:22:@4616.4]
  wire [31:0] core_io_dmem_resp_data; // @[rvtile.scala 30:22:@4616.4]
  wire  core_io_dmem_resp_valid; // @[rvtile.scala 30:22:@4616.4]
  wire [4:0] core_io_ddpath_addr; // @[rvtile.scala 30:22:@4616.4]
  wire [31:0] core_io_ddpath_wdata; // @[rvtile.scala 30:22:@4616.4]
  wire  core_io_ddpath_valid; // @[rvtile.scala 30:22:@4616.4]
  wire [31:0] core_io_ddpath_rdata; // @[rvtile.scala 30:22:@4616.4]
  wire  memarb_clock; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_reset; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_inst_port_req_addr; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_inst_port_req_valid; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_inst_port_resp_data; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_inst_port_resp_valid; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_data_port_req_addr; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_data_port_req_data; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_data_port_req_mfunc; // @[rvtile.scala 32:24:@4619.4]
  wire [1:0] memarb_io_data_port_req_mtype; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_data_port_req_valid; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_data_port_req_ready; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_data_port_resp_data; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_data_port_resp_valid; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_dm_port_req_addr; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_dm_port_req_data; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_dm_port_req_mfunc; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_dm_port_req_valid; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_dm_port_req_ready; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_dm_port_resp_data; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_dm_port_resp_valid; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_waen; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_wden; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_ext_mem_waddr; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_ext_mem_wdata; // @[rvtile.scala 32:24:@4619.4]
  wire [3:0] memarb_io_ext_mem_wmask; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_wardy; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_wdrdy; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_wbvld; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_raen; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_rden; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_ext_mem_raddr; // @[rvtile.scala 32:24:@4619.4]
  wire [31:0] memarb_io_ext_mem_rdata; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_rardy; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_rdrdy; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_clock; // @[rvtile.scala 32:24:@4619.4]
  wire  memarb_io_ext_mem_reset; // @[rvtile.scala 32:24:@4619.4]
  wire  _T_65; // @[rvtile.scala 54:27:@4678.4]
  rvdm dm ( // @[rvtile.scala 29:20:@4613.4]
    .clock(dm_clock),
    .reset(dm_reset),
    .io_dmi_req_bits_op(dm_io_dmi_req_bits_op),
    .io_dmi_req_bits_addr(dm_io_dmi_req_bits_addr),
    .io_dmi_req_bits_data(dm_io_dmi_req_bits_data),
    .io_dmi_req_valid(dm_io_dmi_req_valid),
    .io_dmi_req_ready(dm_io_dmi_req_ready),
    .io_dmi_resp_bits_resp(dm_io_dmi_resp_bits_resp),
    .io_dmi_resp_bits_data(dm_io_dmi_resp_bits_data),
    .io_dmi_resp_valid(dm_io_dmi_resp_valid),
    .io_ddpath_addr(dm_io_ddpath_addr),
    .io_ddpath_wdata(dm_io_ddpath_wdata),
    .io_ddpath_valid(dm_io_ddpath_valid),
    .io_ddpath_rdata(dm_io_ddpath_rdata),
    .io_ddmem_req_addr(dm_io_ddmem_req_addr),
    .io_ddmem_req_data(dm_io_ddmem_req_data),
    .io_ddmem_req_mfunc(dm_io_ddmem_req_mfunc),
    .io_ddmem_req_valid(dm_io_ddmem_req_valid),
    .io_ddmem_req_ready(dm_io_ddmem_req_ready),
    .io_ddmem_resp_data(dm_io_ddmem_resp_data),
    .io_ddmem_resp_valid(dm_io_ddmem_resp_valid),
    .io_rstcore(dm_io_rstcore)
  );
  rvcore core ( // @[rvtile.scala 30:22:@4616.4]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_req_addr(core_io_imem_req_addr),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_resp_data(core_io_imem_resp_data),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_dmem_req_addr(core_io_dmem_req_addr),
    .io_dmem_req_data(core_io_dmem_req_data),
    .io_dmem_req_mfunc(core_io_dmem_req_mfunc),
    .io_dmem_req_mtype(core_io_dmem_req_mtype),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_resp_data(core_io_dmem_resp_data),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_ddpath_addr(core_io_ddpath_addr),
    .io_ddpath_wdata(core_io_ddpath_wdata),
    .io_ddpath_valid(core_io_ddpath_valid),
    .io_ddpath_rdata(core_io_ddpath_rdata)
  );
  rvmemarb memarb ( // @[rvtile.scala 32:24:@4619.4]
    .clock(memarb_clock),
    .reset(memarb_reset),
    .io_inst_port_req_addr(memarb_io_inst_port_req_addr),
    .io_inst_port_req_valid(memarb_io_inst_port_req_valid),
    .io_inst_port_resp_data(memarb_io_inst_port_resp_data),
    .io_inst_port_resp_valid(memarb_io_inst_port_resp_valid),
    .io_data_port_req_addr(memarb_io_data_port_req_addr),
    .io_data_port_req_data(memarb_io_data_port_req_data),
    .io_data_port_req_mfunc(memarb_io_data_port_req_mfunc),
    .io_data_port_req_mtype(memarb_io_data_port_req_mtype),
    .io_data_port_req_valid(memarb_io_data_port_req_valid),
    .io_data_port_req_ready(memarb_io_data_port_req_ready),
    .io_data_port_resp_data(memarb_io_data_port_resp_data),
    .io_data_port_resp_valid(memarb_io_data_port_resp_valid),
    .io_dm_port_req_addr(memarb_io_dm_port_req_addr),
    .io_dm_port_req_data(memarb_io_dm_port_req_data),
    .io_dm_port_req_mfunc(memarb_io_dm_port_req_mfunc),
    .io_dm_port_req_valid(memarb_io_dm_port_req_valid),
    .io_dm_port_req_ready(memarb_io_dm_port_req_ready),
    .io_dm_port_resp_data(memarb_io_dm_port_resp_data),
    .io_dm_port_resp_valid(memarb_io_dm_port_resp_valid),
    .io_ext_mem_waen(memarb_io_ext_mem_waen),
    .io_ext_mem_wden(memarb_io_ext_mem_wden),
    .io_ext_mem_waddr(memarb_io_ext_mem_waddr),
    .io_ext_mem_wdata(memarb_io_ext_mem_wdata),
    .io_ext_mem_wmask(memarb_io_ext_mem_wmask),
    .io_ext_mem_wardy(memarb_io_ext_mem_wardy),
    .io_ext_mem_wdrdy(memarb_io_ext_mem_wdrdy),
    .io_ext_mem_wbvld(memarb_io_ext_mem_wbvld),
    .io_ext_mem_raen(memarb_io_ext_mem_raen),
    .io_ext_mem_rden(memarb_io_ext_mem_rden),
    .io_ext_mem_raddr(memarb_io_ext_mem_raddr),
    .io_ext_mem_rdata(memarb_io_ext_mem_rdata),
    .io_ext_mem_rardy(memarb_io_ext_mem_rardy),
    .io_ext_mem_rdrdy(memarb_io_ext_mem_rdrdy),
    .io_ext_mem_clock(memarb_io_ext_mem_clock),
    .io_ext_mem_reset(memarb_io_ext_mem_reset)
  );
  assign _T_65 = dm_io_rstcore | reset; // @[rvtile.scala 54:27:@4678.4]
  assign io_dmi_req_ready = dm_io_dmi_req_ready;
  assign io_dmi_resp_bits_resp = dm_io_dmi_resp_bits_resp;
  assign io_dmi_resp_bits_data = dm_io_dmi_resp_bits_data;
  assign io_dmi_resp_valid = dm_io_dmi_resp_valid;
  assign io_ext_mem_waen = memarb_io_ext_mem_waen;
  assign io_ext_mem_wden = memarb_io_ext_mem_wden;
  assign io_ext_mem_waddr = memarb_io_ext_mem_waddr;
  assign io_ext_mem_wdata = memarb_io_ext_mem_wdata;
  assign io_ext_mem_wmask = memarb_io_ext_mem_wmask;
  assign io_ext_mem_raen = memarb_io_ext_mem_raen;
  assign io_ext_mem_rden = memarb_io_ext_mem_rden;
  assign io_ext_mem_raddr = memarb_io_ext_mem_raddr;
  assign io_ext_mem_clock = memarb_io_ext_mem_clock;
  assign io_ext_mem_reset = memarb_io_ext_mem_reset;
  assign dm_clock = clock;
  assign dm_reset = reset;
  assign dm_io_dmi_req_bits_op = io_dmi_req_bits_op;
  assign dm_io_dmi_req_bits_addr = io_dmi_req_bits_addr;
  assign dm_io_dmi_req_bits_data = io_dmi_req_bits_data;
  assign dm_io_dmi_req_valid = io_dmi_req_valid;
  assign dm_io_ddpath_rdata = core_io_ddpath_rdata;
  assign dm_io_ddmem_req_ready = memarb_io_dm_port_req_ready;
  assign dm_io_ddmem_resp_data = memarb_io_dm_port_resp_data;
  assign dm_io_ddmem_resp_valid = memarb_io_dm_port_resp_valid;
  assign core_clock = clock;
  assign core_reset = _T_65;
  assign core_io_imem_resp_data = memarb_io_inst_port_resp_data;
  assign core_io_imem_resp_valid = memarb_io_inst_port_resp_valid;
  assign core_io_dmem_req_ready = memarb_io_data_port_req_ready;
  assign core_io_dmem_resp_data = memarb_io_data_port_resp_data;
  assign core_io_dmem_resp_valid = memarb_io_data_port_resp_valid;
  assign core_io_ddpath_addr = dm_io_ddpath_addr;
  assign core_io_ddpath_wdata = dm_io_ddpath_wdata;
  assign core_io_ddpath_valid = dm_io_ddpath_valid;
  assign memarb_clock = clock;
  assign memarb_reset = reset;
  assign memarb_io_inst_port_req_addr = core_io_imem_req_addr;
  assign memarb_io_inst_port_req_valid = core_io_imem_req_valid;
  assign memarb_io_data_port_req_addr = core_io_dmem_req_addr;
  assign memarb_io_data_port_req_data = core_io_dmem_req_data;
  assign memarb_io_data_port_req_mfunc = core_io_dmem_req_mfunc;
  assign memarb_io_data_port_req_mtype = core_io_dmem_req_mtype;
  assign memarb_io_data_port_req_valid = core_io_dmem_req_valid;
  assign memarb_io_dm_port_req_addr = dm_io_ddmem_req_addr;
  assign memarb_io_dm_port_req_data = dm_io_ddmem_req_data;
  assign memarb_io_dm_port_req_mfunc = dm_io_ddmem_req_mfunc;
  assign memarb_io_dm_port_req_valid = dm_io_ddmem_req_valid;
  assign memarb_io_ext_mem_wardy = io_ext_mem_wardy;
  assign memarb_io_ext_mem_wdrdy = io_ext_mem_wdrdy;
  assign memarb_io_ext_mem_wbvld = io_ext_mem_wbvld;
  assign memarb_io_ext_mem_rdata = io_ext_mem_rdata;
  assign memarb_io_ext_mem_rardy = io_ext_mem_rardy;
  assign memarb_io_ext_mem_rdrdy = io_ext_mem_rdrdy;
endmodule
module rv32i_fpga( // @[:@4681.2]
  input         clock, // @[:@4682.4]
  input         reset, // @[:@4683.4]
  input  [1:0]  io_dmi_req_bits_op, // @[:@4684.4]
  input  [6:0]  io_dmi_req_bits_addr, // @[:@4684.4]
  input  [31:0] io_dmi_req_bits_data, // @[:@4684.4]
  input         io_dmi_req_valid, // @[:@4684.4]
  output        io_dmi_req_ready, // @[:@4684.4]
  output [1:0]  io_dmi_resp_bits_resp, // @[:@4684.4]
  output [31:0] io_dmi_resp_bits_data, // @[:@4684.4]
  output        io_dmi_resp_valid, // @[:@4684.4]
  input         io_dmi_resp_ready, // @[:@4684.4]
  output        io_ext_mem_waen, // @[:@4684.4]
  output        io_ext_mem_wden, // @[:@4684.4]
  output [31:0] io_ext_mem_waddr, // @[:@4684.4]
  output [31:0] io_ext_mem_wdata, // @[:@4684.4]
  output [3:0]  io_ext_mem_wmask, // @[:@4684.4]
  input         io_ext_mem_wardy, // @[:@4684.4]
  input         io_ext_mem_wdrdy, // @[:@4684.4]
  input         io_ext_mem_wbvld, // @[:@4684.4]
  output        io_ext_mem_raen, // @[:@4684.4]
  output        io_ext_mem_rden, // @[:@4684.4]
  output [31:0] io_ext_mem_raddr, // @[:@4684.4]
  input  [31:0] io_ext_mem_rdata, // @[:@4684.4]
  input         io_ext_mem_rardy, // @[:@4684.4]
  input         io_ext_mem_rdrdy, // @[:@4684.4]
  output        io_ext_mem_clock, // @[:@4684.4]
  output        io_ext_mem_reset // @[:@4684.4]
);
  wire  rvtile_clock; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_reset; // @[rvfpga.scala 24:24:@4686.4]
  wire [1:0] rvtile_io_dmi_req_bits_op; // @[rvfpga.scala 24:24:@4686.4]
  wire [6:0] rvtile_io_dmi_req_bits_addr; // @[rvfpga.scala 24:24:@4686.4]
  wire [31:0] rvtile_io_dmi_req_bits_data; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_dmi_req_valid; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_dmi_req_ready; // @[rvfpga.scala 24:24:@4686.4]
  wire [1:0] rvtile_io_dmi_resp_bits_resp; // @[rvfpga.scala 24:24:@4686.4]
  wire [31:0] rvtile_io_dmi_resp_bits_data; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_dmi_resp_valid; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_waen; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_wden; // @[rvfpga.scala 24:24:@4686.4]
  wire [31:0] rvtile_io_ext_mem_waddr; // @[rvfpga.scala 24:24:@4686.4]
  wire [31:0] rvtile_io_ext_mem_wdata; // @[rvfpga.scala 24:24:@4686.4]
  wire [3:0] rvtile_io_ext_mem_wmask; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_wardy; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_wdrdy; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_wbvld; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_raen; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_rden; // @[rvfpga.scala 24:24:@4686.4]
  wire [31:0] rvtile_io_ext_mem_raddr; // @[rvfpga.scala 24:24:@4686.4]
  wire [31:0] rvtile_io_ext_mem_rdata; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_rardy; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_rdrdy; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_clock; // @[rvfpga.scala 24:24:@4686.4]
  wire  rvtile_io_ext_mem_reset; // @[rvfpga.scala 24:24:@4686.4]
  rvtile rvtile ( // @[rvfpga.scala 24:24:@4686.4]
    .clock(rvtile_clock),
    .reset(rvtile_reset),
    .io_dmi_req_bits_op(rvtile_io_dmi_req_bits_op),
    .io_dmi_req_bits_addr(rvtile_io_dmi_req_bits_addr),
    .io_dmi_req_bits_data(rvtile_io_dmi_req_bits_data),
    .io_dmi_req_valid(rvtile_io_dmi_req_valid),
    .io_dmi_req_ready(rvtile_io_dmi_req_ready),
    .io_dmi_resp_bits_resp(rvtile_io_dmi_resp_bits_resp),
    .io_dmi_resp_bits_data(rvtile_io_dmi_resp_bits_data),
    .io_dmi_resp_valid(rvtile_io_dmi_resp_valid),
    .io_ext_mem_waen(rvtile_io_ext_mem_waen),
    .io_ext_mem_wden(rvtile_io_ext_mem_wden),
    .io_ext_mem_waddr(rvtile_io_ext_mem_waddr),
    .io_ext_mem_wdata(rvtile_io_ext_mem_wdata),
    .io_ext_mem_wmask(rvtile_io_ext_mem_wmask),
    .io_ext_mem_wardy(rvtile_io_ext_mem_wardy),
    .io_ext_mem_wdrdy(rvtile_io_ext_mem_wdrdy),
    .io_ext_mem_wbvld(rvtile_io_ext_mem_wbvld),
    .io_ext_mem_raen(rvtile_io_ext_mem_raen),
    .io_ext_mem_rden(rvtile_io_ext_mem_rden),
    .io_ext_mem_raddr(rvtile_io_ext_mem_raddr),
    .io_ext_mem_rdata(rvtile_io_ext_mem_rdata),
    .io_ext_mem_rardy(rvtile_io_ext_mem_rardy),
    .io_ext_mem_rdrdy(rvtile_io_ext_mem_rdrdy),
    .io_ext_mem_clock(rvtile_io_ext_mem_clock),
    .io_ext_mem_reset(rvtile_io_ext_mem_reset)
  );
  assign io_dmi_req_ready = rvtile_io_dmi_req_ready;
  assign io_dmi_resp_bits_resp = rvtile_io_dmi_resp_bits_resp;
  assign io_dmi_resp_bits_data = rvtile_io_dmi_resp_bits_data;
  assign io_dmi_resp_valid = rvtile_io_dmi_resp_valid;
  assign io_ext_mem_waen = rvtile_io_ext_mem_waen;
  assign io_ext_mem_wden = rvtile_io_ext_mem_wden;
  assign io_ext_mem_waddr = rvtile_io_ext_mem_waddr;
  assign io_ext_mem_wdata = rvtile_io_ext_mem_wdata;
  assign io_ext_mem_wmask = rvtile_io_ext_mem_wmask;
  assign io_ext_mem_raen = rvtile_io_ext_mem_raen;
  assign io_ext_mem_rden = rvtile_io_ext_mem_rden;
  assign io_ext_mem_raddr = rvtile_io_ext_mem_raddr;
  assign io_ext_mem_clock = rvtile_io_ext_mem_clock;
  assign io_ext_mem_reset = rvtile_io_ext_mem_reset;
  assign rvtile_clock = clock;
  assign rvtile_reset = reset;
  assign rvtile_io_dmi_req_bits_op = io_dmi_req_bits_op;
  assign rvtile_io_dmi_req_bits_addr = io_dmi_req_bits_addr;
  assign rvtile_io_dmi_req_bits_data = io_dmi_req_bits_data;
  assign rvtile_io_dmi_req_valid = io_dmi_req_valid;
  assign rvtile_io_ext_mem_wardy = io_ext_mem_wardy;
  assign rvtile_io_ext_mem_wdrdy = io_ext_mem_wdrdy;
  assign rvtile_io_ext_mem_wbvld = io_ext_mem_wbvld;
  assign rvtile_io_ext_mem_rdata = io_ext_mem_rdata;
  assign rvtile_io_ext_mem_rardy = io_ext_mem_rardy;
  assign rvtile_io_ext_mem_rdrdy = io_ext_mem_rdrdy;
endmodule
